`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "XILINX"
`pragma protect encrypt_agent_info = "Xilinx Encryption Tool 2020.2"
`pragma protect key_keyowner = "Cadence Design Systems.", key_keyname = "cds_rsa_key", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`pragma protect key_block
C0oJF2SuMa6l5UTKL3oQ8NzIzSt0InrgoMNkISrJfbH+L4MIoyjcJGHLfWlSoL8sgNnJJnewfJpv
YfYxDbNsYw==

`pragma protect key_keyowner = "Synopsys", key_keyname = "SNPS-VCS-RSA-2", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`pragma protect key_block
T73gREUbEeEcadgcm0Fok6jWAkVLLIAj0g8M1ElpcxW4VzJb7Eg2z1clk1vvjr+ennzWkPDdCqSR
7g1wInRiACjYhCUiSW+M3ZYhyRrZqbojKW6+M6XtNNyn9fcoc4CNqjb1z0dKzQN2Ed5VjTvH1b3k
XUlVT3178PUueN/MvG8=

`pragma protect key_keyowner = "Aldec", key_keyname = "ALDEC15_001", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`pragma protect key_block
Zp3QCPiy/URa5u3qn57TB9bhSAk9uQ0biVaxe4uWXuJ7pemvtklJ69FjvHdb5FlPJdQntbtpj0/f
edX5k/wcAwuTS7H7DPI0Ws1Bqz6CKOD4xaTHv2oslshZRaRQvIrmdN4Rw/5qp2ZSG06Xi1hSxVvK
Jg0eu8PcJGqYXLYgb5QC7INxxreeqds+4xrIlpd1HK3jxui3Whj9er/dQnJZ+TMX0wEAQBixOsBG
gnogY/28/lCm/qKY5uKuvCtCyYlW7kpiaqwLtVfSOPUBakWeQunH87r+ZPutRUEJSHSqQNJG7+4t
N3FqL8iQR3HwsFNLhMXnNGbvWTOug7VJ8JNqTQ==

`pragma protect key_keyowner = "ATRENTA", key_keyname = "ATR-SG-2015-RSA-3", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`pragma protect key_block
WlpHIH6+59sUqAlQSWev+VnSCbtuwXM7bkHr4rCUbCJtTzC2OvCApSZHHGXFjCeg/5bXtIcJ+Z6g
fgSBcRGjcyg06GJjida88LkRfX1zal7u1LQZ/b6AKUY6GJXA8fgPa16oGYoXZCRglkTA0usTHpvU
7zVrw1GSAcV1Rqk2JMMs/7odJmb3bPnHsmAPM7GmZmff/DMbNQTrS2NWKvl6Y68UbMLeI/+wL6n/
tED2pvdOQm6tYXELI+YSUhIVfyK/Rcy3S1S8Nqa8E/034z15I/GKyVdJpVb6rX0V+sIfvzBHjNBp
v5XcsEe+J5UR6CR5b+OuhKT8AVnqMVmm2lrdHQ==

`pragma protect key_keyowner = "Mentor Graphics Corporation", key_keyname = "MGC-VELOCE-RSA", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`pragma protect key_block
s1auGT8s07pA5X1CC1iqJE3xKUF37HebCmECcARl84x+0IqQT4kdboNEDw+7/H6a6MdaMRGhTeef
X922orJDDURsbC8Xt2TrwldYajGk8jNMzNqfIuVWMLvijNTGfyPl4kUyXOri6Y/HpCMAiqQTUn/0
C7m1aWIFJDiPm2SuNr8=

`pragma protect key_keyowner = "Mentor Graphics Corporation", key_keyname = "MGC-VERIF-SIM-RSA-2", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`pragma protect key_block
Ei7FxD+k4QZBqit678M6N0vzExc2reWl5rdBjfOMq2fMZ/ljOAmwMn+uaUXPYEQMXm+/5admVo2G
/C2zPOsusl+osaeETBe+bh8KF27lPvYzGK4ziQR3Hi3I30oOyo4V9GjRSEZz7reDE2SNeUnB8RVz
B3g93eF5IwwjnW2AwNtgf6E4gvYQeRoPk9UAN0duY/fH60P0Wx3FUEcN5sey/ExJ3MmU7VCZH9/v
U/6Wj0BdwAleZFNFfBxNyQHnVS/wE35qsyb1cOonZu/fsEMcbav/p03XIvoRmdl0X5cZt8RcQdav
ojYJeAb/sCrZOqzm0FpR5M4Owh4aRCCj/kNbrw==

`pragma protect key_keyowner = "Real Intent", key_keyname = "RI-RSA-KEY-1", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`pragma protect key_block
wY9QtmtV84Now9Kq9cA7AwRQ7O4mNcEX8FDE3uCBJzno/JF7N3J321QnQ0dxXW/iXhyYnlCuC2Va
oOnDA5SidFCVZ9Q7gmc5vUg0fph8Wng5BwwPJ8XUP1mHqYKHs8vYtA9G4lSTuUBj9jRhLQQkf3TV
IE1yzmILHl/aUpBqmkjJ6mRZo8dQS2i4Yc9NH6BTPRQDS0yFgh8/mexim1nT6vgTgNf14h7omDPI
amNp3Aafutw6k/xU8eqYRWR7pytlYHCia7+HHjwBI7dUl7T4UjmG1q3x87TmcZ1q2u9vHJsEIMMV
34EVPExsKjtifd6Dd5mguDr8rIKSaRCF2tjtkw==

`pragma protect key_keyowner = "Metrics Technologies Inc.", key_keyname = "DSim", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`pragma protect key_block
eVM+E5yFaaEW0df0uVjFsuziATF5vfG4cSmmBEuGSLcO7WzDsopPqRvwLQ/P2P+nqdPLXPj7At7t
U0/Uoeb8h2mikT0Y3O4xYwsot79/uJ/fh4wLf0kCYLBvH8+4eGdt+OZbMATC8w3MMDU/Ztey+dWx
VXf8/lyxU6R/Y2RF1AU6lGpB/rar5mImrHV90febD3ItbvH1TmTnj8NJDMO8jvm4xuUtJojg0Nmj
43DvyUbmQCOK+8gCjCOyQhPMdTh5p+mx8x6fIuHL935kMkcogRtUZp/3Xp6dlMP35OJpsEogX209
xaOi6daJVsalpJOhvKwOEwRsC1uQD7w/BNt/KQ==

`pragma protect key_keyowner = "Xilinx", key_keyname = "xilinxt_2020_08", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`pragma protect key_block
RPpz5aiA1FU3P+Y4nj5b2duqFntW7YLQveNMMRIIbWzptbnClOymdlEWJll+G1/aDsYWhqtwulkx
/ZfVvXbuYhuDIgOmOQTYxBkrYPxDN9SIGBuyZAN8s9OShmCUJ5cNv+nog+9fJ6Bvh3UTbZ2IPT7Q
I4tpfDJnw8MlFrTEULEYa4JuAe4NHW9lwZI9FVlNY/53wP8EYxF8OJmPPts7wQSzH7XnVytpXV+p
wZ4L0VtXEvZSCC+7AAftazTSHzxX2p6FbWl55UOIHXC+rxevOa+eATCnR8PO0GwNB5VyH6IhvH04
f4ifslvamlFYShLgBLBEOjfwmCe/0MdAwDeQ7A==

`pragma protect data_method = "AES128-CBC"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 3136)
`pragma protect data_block
SqC3s74hTjR+1MFnTJCcueRiGlzqJFhYh6eWPKALuL7KYy2lbYdsr/9zqMa/25XHfuvUp4fSvxcF
eSSe5S8ZPx7owrOIEftAknToJrUrCvGFaksghVnGqwI3ZfU/sUDnAK6bhJQNz6FcAYODJ1ro33/s
IcKifDukxb4Fk/vPWLjGodiyLe/sE39sZJgHrSNbsRp95OG3EFTvxqQBtdgn8tWbNqJKARxMispc
fwF8CXBGGM/T6aA84rQxP1OrDzGE/H5Vkb4FeKx3NOvWzTA5aMsSv1I6Af3WFQ0g9e51henrX2Ql
P1USthNS06xut2D0wh3RIn3ZhnWDnTbya4tFFCf73tBGj4ju1l9i6uFAEMCFbuoa7gQogyzj+Xpy
PGu0fxBMKqmIM+488Ghq3iM6HC/JYmOxKU1yMlBVD0FTKUAm+vnD8YF4bQOn+cOOv+8iGsluCEEb
sI1acyCsQ0ANhccB14q1kfKyKCLDU/Q/WfKKERSGMfITaQC/97G7RZgDs6SS5VLlukKlbrb5J5N3
5fqrp227qNGzkORjIuIRbN+iJCTv3J5paswGpvq2p7CWb8gs7Bs6MsqQAFrUpnLD4ULvoZ2R6Y3h
NmcjtM3BWBIwjIcZRvKW71wZY9mIe9zHlUS/KXl9ABqWycGuKjn4IE6tE01qFhvy6RcosOExn3sY
uzRk4HBEAFw5rODNOSaabn96bq1Rq1gEkQOdyFChPHn6HDkLBD6YcFB6Fatk8GP2v/V4cB7jQQJN
2vgk41xzvX79CDu1SIiWkdoUtT5CXrXEvqkQNPnhIHLEf69LhXv2Tg7EszxeYOXZikgAJSwJ6KiF
PV9zKR20oUSoxB6eGJFmTZmLrITCAw8AXIGy1Kob1/oGEE0/6Hlp+wb/ULpAscIaGZ9kSCfOaFQc
EOV3EbROJ9JG7a2FPvvsyqs6923GZ/352facXpFjmVlr3L4CkKHTAkQTZ21JMTgG2s6VdlmyGBLM
hcCXBa0MgsPbau2rqkZYhwOnBmWWpeFMnV51TGK+9DdfiDUibVzTtbEGB1nn+6IdGb2fvOceKpw0
qlO1z4ol7vB0ZdAIwNCehSfq9awhe7iune/YeGQNRSjCvoVrh/GIk5YQ5DzunhOLy0KS2JHd5mD/
znZZ3n9y3FyM2jykTIrK/OX2/ezyDXcL4ASmcR3WS4fn1DTBGwIwynYu2CB94X2elBMiWiQJ7Dkx
w+CPHemf8eOKEKD9Dgm7iIpCS+qkj+u+ArSvrGFZdRi0F2IdrvdISAKBvvrG0mTpijQWtg3/ZEzG
00lTMIgEbRqis9TKeL9HRT9KDu8nRNt4P+oTTiJvl5/QGA3QU1eVpPPuLoobpRSoyFSwQV7OnJsB
eTexBHuXnsf/gtepaEI7YJVjliwzUQa18Sq/P5CRvBkAGfqugmTDhMZR3tRpVTSbQSTAABeqN/LG
iuzit6yaoThzmGd8LzvBh+bx1+6oHre+lWy9Wi3QdYXlBvnBY4DwiGzQXX1bcu3KEThfPZcihiS3
ZYnVR5CigMFXAWXwpwfKiqmL5LRgW72qIFbYUDMQjau48EI42y1BW7RhkkAy5EWlBtyWlS7NBkYv
anEI+iUblt3Uk2rw06G1FNVlthEKQg3Nz6FJWEa2vnoK8YcN8Tejsq8CqUCFYeGzmNOmHEsm3JQ2
SO15xx1XCZlA6zFPxeFr2DVw1dxrASK/3n0fRvXhdFlEC3fAKbKUEg0w8NGB0+7BQ63UVGnybTtm
VJHvZekZSOKI++MI+Z0zM2Xrc/NIWAWsE5B5jY1ANZkWGRBi4bdqPHHmFtI1gui0oiXhbiSCDIJ7
eCEyyHs/ZPyf7tnAt4mjaI+6JU1FXrF8SFrBq4fbqFcijDXik/kcZreYaxZaJcZjD5pA3JLxC97D
NoSCDk0xMHUN9pIf0Q/R3d+nY5bQSDefRz7a7Szg0B6ual1fEEe2Tity9ncGWLl6aOflebTx7mnH
ZiktbG9iW4dIe+vxWQhtH+cqf1xR3OzSO//jZhNsP5dPpx4AuCj/IPqbYRkh6FdEe2jFjJOOEeoB
XR8FMjoe7AW5BJd6FqergOrOSgmA5NMeGbf2PNdFgd4nqzx4etHv+fL6NKBkdvwNKr3iASKA9ZHq
vtm0THi7VaKRhzABGjmGsx/mqYVzep7uMyGfLb2XvjVuNFoqm9GX6uoc9TS+Dg5Y4oCtK8Mna1Kp
Hf58KoRST7jwnglSUuoxFT3P7RbjfRKqwegD+J7fkzyv76Yrjrw+oFufT35Qtrq/6sCiY0fp9lVJ
Iu2TA+vDtyAj6Uk+pJ2TQ/qvqzQrm7y/IYKNFHxqiwNlTMJ1bmBdw0ipdORNHmpWgVj4QeUm/8nx
zO/HSabzVysPV3ApmWBd/+RV2ZMSASmN7ruOE6U7siDTJuOaBNMOS/7Z2CkvcGLFxuiibN+H67/q
RkcU+jNAFM9SCQulFmC/deWO+jkVNFRUuQmsA0YQ9XAUF8azZvVkARrJmzNaTeak06XY3mEGzPtC
WMw77q+cKImqHrm3fXz2RqQPaGZqzxeQelirPMiVcsohzI1cj84s/S4zLd+3U7pnS5nw9mYfOc9g
woyBePuT83oIz+3siZowRlm9qUd6z7lT6yM0s0kNtU/3mcaArX7GnOcrEd6ku2/+aH9Xem2qKEH4
qoxBE5Riqvdhlj9VfJtO4S8rBqr8fN076Ti5XIgysv5uTmEuQ9naakNspDwk30h5k4sIh7YiNUF5
Xzy1Srm90LmE2GJRNlzC9Xp78qYXVJq7RIRVSQxh/7CS0bADR0rtnYA+2YTI4ISd1BlNNNSiIdGb
I9tPTrgXzidaJOp7TSbv7kZ2Jbm83Pd4lp63ur4KzjflbPuJj3mrFPYphRK4oJb41EndgJcKWSFY
IGQlg2b0PwqCZn1eDxSRe1Y86vaxclrnCioDjNiGQ/kI85mMNs4KfvMc7BNcwdHdIIQT87bR15Yb
S7jotQLwWN3kBD97dSNDmQSLihXsDyxHBZtHKwrmcbhMbSPE4RZtVWsBxOPrPcUfKh6vIE3gT+ja
Cu5D5g22clkdt47GkBUm3d9GAM4BK6Cfc+2p+u2Nhkaok/QjGiUNIPdCOybKKoSkhTWKnTnVIDmg
IkuM/7NteTgk7CXhHkhXANjg+81MpP8TeII3c95gAvPOrE22fKmfHGmDHg0GRHhm1iCpGGFSu3bo
JBrt5M1Z8M7IYtoVlPJDhBHYfUBqN0caoLcSOC5WRcniYNm51EP8xkBXm1tJpCuZLrWwgyJM7dpn
syhR9Jp3k13YRk5Jde4TyuYwUlKr58iARig7FZDzqP8h+FiGJWgePxDVHHY6EfWPXZVGG6QcGVYu
3mzzc8AvNCD7gh4cIrA1EZpGABmpKjBQU8ARWz4wrwiCanjBQWen8jK+CknG5ChTgg9N/676+SvS
ZryppMwbmCbA54toKq6G+fFxawCNdS0BwD9BN1Y6P7kvI6cYixdQd4WUm+j6HpqXI4sXJ8z+vt/T
ZeW9fhLhx9MGbRoRjtTAdD7nB6puLBMGVqQ8ac0Z+oENbwV0ctdFciLDxZN/4bU73p9qxyJeC5p3
1DqV8+Ryu5jk06S2IExsrui+mTi/bFpWvO4Z93Oa4lW+3Rp4Es0PdpMQT0eqFPxz5BGkGEnXYEgR
FqxQspiCgntRY7V+BW4e2ok3oFZ64ZEQnDoeK7j9kmu1JBhJ2bYBg2cVVDA94JOVji4Zcp8k3Iek
fZaSBl/vg9ekpzShzGVeP4RAvoA7aL9YVcCR5r1lhetT3gF5KLI+e/JocxA8duA5LqbZtDXHmQp9
DGzAKbzcru1uY9KOz+s8O7LLGY7579cjlFb+WmXb/87RUR48jl/r5Kxt1AIO4ZOaQZKaqwPRXhVW
gxV2wQSeWtYztuZVlYsnTuaSUHmryYGB+K/VXVdsrfF+VB4ZPYCfASm8EQz7j/KvEEN/jRqDWio5
o2Q2W3JXLs9UC8Uo+jcEuPTWWkQSrMWC+BQ/Pf4+d61aOqOn8jH7MreGgdaKCUFqLxvwWafjNLaA
wsrac5ntcq/qjUcH+5ehN928cCZbhKf+Kbjf8gZNXQudwbNTajX1Kw6D9i5CreX2g0zZoYsDqs/w
5JPwM2OT7To3BliMYR3FE73cWVk8AeUiG7Ad47lckLPHbvBVHqrRwZf+DBNUSk0/9S2ccLMR4/ah
ow==
`pragma protect end_protected
