`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "XILINX"
`pragma protect encrypt_agent_info = "Xilinx Encryption Tool 2020.2"
`pragma protect key_keyowner = "Cadence Design Systems.", key_keyname = "cds_rsa_key", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`pragma protect key_block
C0oJF2SuMa6l5UTKL3oQ8NzIzSt0InrgoMNkISrJfbH+L4MIoyjcJGHLfWlSoL8sgNnJJnewfJpv
YfYxDbNsYw==

`pragma protect key_keyowner = "Synopsys", key_keyname = "SNPS-VCS-RSA-2", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`pragma protect key_block
T73gREUbEeEcadgcm0Fok6jWAkVLLIAj0g8M1ElpcxW4VzJb7Eg2z1clk1vvjr+ennzWkPDdCqSR
7g1wInRiACjYhCUiSW+M3ZYhyRrZqbojKW6+M6XtNNyn9fcoc4CNqjb1z0dKzQN2Ed5VjTvH1b3k
XUlVT3178PUueN/MvG8=

`pragma protect key_keyowner = "Aldec", key_keyname = "ALDEC15_001", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`pragma protect key_block
Zp3QCPiy/URa5u3qn57TB9bhSAk9uQ0biVaxe4uWXuJ7pemvtklJ69FjvHdb5FlPJdQntbtpj0/f
edX5k/wcAwuTS7H7DPI0Ws1Bqz6CKOD4xaTHv2oslshZRaRQvIrmdN4Rw/5qp2ZSG06Xi1hSxVvK
Jg0eu8PcJGqYXLYgb5QC7INxxreeqds+4xrIlpd1HK3jxui3Whj9er/dQnJZ+TMX0wEAQBixOsBG
gnogY/28/lCm/qKY5uKuvCtCyYlW7kpiaqwLtVfSOPUBakWeQunH87r+ZPutRUEJSHSqQNJG7+4t
N3FqL8iQR3HwsFNLhMXnNGbvWTOug7VJ8JNqTQ==

`pragma protect key_keyowner = "ATRENTA", key_keyname = "ATR-SG-2015-RSA-3", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`pragma protect key_block
WlpHIH6+59sUqAlQSWev+VnSCbtuwXM7bkHr4rCUbCJtTzC2OvCApSZHHGXFjCeg/5bXtIcJ+Z6g
fgSBcRGjcyg06GJjida88LkRfX1zal7u1LQZ/b6AKUY6GJXA8fgPa16oGYoXZCRglkTA0usTHpvU
7zVrw1GSAcV1Rqk2JMMs/7odJmb3bPnHsmAPM7GmZmff/DMbNQTrS2NWKvl6Y68UbMLeI/+wL6n/
tED2pvdOQm6tYXELI+YSUhIVfyK/Rcy3S1S8Nqa8E/034z15I/GKyVdJpVb6rX0V+sIfvzBHjNBp
v5XcsEe+J5UR6CR5b+OuhKT8AVnqMVmm2lrdHQ==

`pragma protect key_keyowner = "Mentor Graphics Corporation", key_keyname = "MGC-VELOCE-RSA", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`pragma protect key_block
s1auGT8s07pA5X1CC1iqJE3xKUF37HebCmECcARl84x+0IqQT4kdboNEDw+7/H6a6MdaMRGhTeef
X922orJDDURsbC8Xt2TrwldYajGk8jNMzNqfIuVWMLvijNTGfyPl4kUyXOri6Y/HpCMAiqQTUn/0
C7m1aWIFJDiPm2SuNr8=

`pragma protect key_keyowner = "Mentor Graphics Corporation", key_keyname = "MGC-VERIF-SIM-RSA-2", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`pragma protect key_block
Ei7FxD+k4QZBqit678M6N0vzExc2reWl5rdBjfOMq2fMZ/ljOAmwMn+uaUXPYEQMXm+/5admVo2G
/C2zPOsusl+osaeETBe+bh8KF27lPvYzGK4ziQR3Hi3I30oOyo4V9GjRSEZz7reDE2SNeUnB8RVz
B3g93eF5IwwjnW2AwNtgf6E4gvYQeRoPk9UAN0duY/fH60P0Wx3FUEcN5sey/ExJ3MmU7VCZH9/v
U/6Wj0BdwAleZFNFfBxNyQHnVS/wE35qsyb1cOonZu/fsEMcbav/p03XIvoRmdl0X5cZt8RcQdav
ojYJeAb/sCrZOqzm0FpR5M4Owh4aRCCj/kNbrw==

`pragma protect key_keyowner = "Real Intent", key_keyname = "RI-RSA-KEY-1", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`pragma protect key_block
wY9QtmtV84Now9Kq9cA7AwRQ7O4mNcEX8FDE3uCBJzno/JF7N3J321QnQ0dxXW/iXhyYnlCuC2Va
oOnDA5SidFCVZ9Q7gmc5vUg0fph8Wng5BwwPJ8XUP1mHqYKHs8vYtA9G4lSTuUBj9jRhLQQkf3TV
IE1yzmILHl/aUpBqmkjJ6mRZo8dQS2i4Yc9NH6BTPRQDS0yFgh8/mexim1nT6vgTgNf14h7omDPI
amNp3Aafutw6k/xU8eqYRWR7pytlYHCia7+HHjwBI7dUl7T4UjmG1q3x87TmcZ1q2u9vHJsEIMMV
34EVPExsKjtifd6Dd5mguDr8rIKSaRCF2tjtkw==

`pragma protect key_keyowner = "Metrics Technologies Inc.", key_keyname = "DSim", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`pragma protect key_block
eVM+E5yFaaEW0df0uVjFsuziATF5vfG4cSmmBEuGSLcO7WzDsopPqRvwLQ/P2P+nqdPLXPj7At7t
U0/Uoeb8h2mikT0Y3O4xYwsot79/uJ/fh4wLf0kCYLBvH8+4eGdt+OZbMATC8w3MMDU/Ztey+dWx
VXf8/lyxU6R/Y2RF1AU6lGpB/rar5mImrHV90febD3ItbvH1TmTnj8NJDMO8jvm4xuUtJojg0Nmj
43DvyUbmQCOK+8gCjCOyQhPMdTh5p+mx8x6fIuHL935kMkcogRtUZp/3Xp6dlMP35OJpsEogX209
xaOi6daJVsalpJOhvKwOEwRsC1uQD7w/BNt/KQ==

`pragma protect key_keyowner = "Xilinx", key_keyname = "xilinxt_2020_08", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`pragma protect key_block
RPpz5aiA1FU3P+Y4nj5b2duqFntW7YLQveNMMRIIbWzptbnClOymdlEWJll+G1/aDsYWhqtwulkx
/ZfVvXbuYhuDIgOmOQTYxBkrYPxDN9SIGBuyZAN8s9OShmCUJ5cNv+nog+9fJ6Bvh3UTbZ2IPT7Q
I4tpfDJnw8MlFrTEULEYa4JuAe4NHW9lwZI9FVlNY/53wP8EYxF8OJmPPts7wQSzH7XnVytpXV+p
wZ4L0VtXEvZSCC+7AAftazTSHzxX2p6FbWl55UOIHXC+rxevOa+eATCnR8PO0GwNB5VyH6IhvH04
f4ifslvamlFYShLgBLBEOjfwmCe/0MdAwDeQ7A==

`pragma protect data_method = "AES128-CBC"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 135968)
`pragma protect data_block
SqC3s74hTjR+1MFnTJCcueRiGlzqJFhYh6eWPKALuL7KYy2lbYdsr/9zqMa/25XHfuvUp4fSvxcF
eSSe5S8ZPx7owrOIEftAknToJrUrCvGMYBsNp3BdTB93XRs1RFWZNtaoSVonGTw+YP5binO4dbaf
VNgcOlubifNVnSvYahQ0980IfJpWD6b5pcOVM2qjEl57R/Abykbs+uMkM/W4rlH0Qp/fSg5Vp2C4
n1AjRdNZgO0GuQxkb1dFLeqOECdGyKHvxqjiW28IG6U131HK7akF8ncKafbvgEKkDhP6kkGavTWS
voyZR6ifx+w/KgR3WQvPYr+R5h0gNFkcAiGgA6iRA39O/ArrGpV75E0nzzaPmVhm7QQ+9sYSGHyu
+7rxcqyKRpQH899Oe8ytCFYZBUUU5LJ5dQOnh3bk4LQxPl12JwjrhwHrGhMQjNOobIsNCQ3T447O
VF0NwpI1RnZL0z/td5Z18Jy+UTSqNkOCouW2l46luAy+REfRaSBDTRXeZI6+j2spdPN1cHuy6wHN
KWtFfbaQuXei6irSX2mevHyrNfKFHAv2zvlINUtnPxy5sKQf0Wqahd6Wfvj94X+0VJ3zkOkcPe20
x9TkjBXPvT5EdBIzDz2WDjnZuSeCKUzGMPDgiN5g4Py1KX4d+2Su7zi7U56b4v4e5beHmKHsvfv7
IwJ+oMAQvPaPlr08MMv/PEfRwY+hrd87it/Mdt0zNgnuNZnxb4zZShyQ8kpzeISpaIGyPyT4ShiG
dYtNtanDlouARjw8DTxaZzHbERnrWlLNS+0JaHPLrHBzMg40QeJ+Lbq8qoHSW9/+QpvV34Cs3np0
ihk81ZWcnjpT4i9lxkHl/mpoKvj6Nr0ms07nqhcitSn0IKSeK0nQ8AixzJOVoE5ANFr0NxIHLSjy
uV4wTjpdyDbYcbZFaLmcuGP8+bZe0DYynd0HsTzfkn7Oie/JX4TxoWZOpsB+RiCvCxLM7ocmsreE
SxI6lFa2UW5HOeuBSqSkj91ZMJv65gQ8iJe/JRsNGv7RDkS/ObJh+USJJ14Ih2WssNjyIX6JhGGC
25F4SAC5hzHogQsAPIqJpAOyL5tqhCwSPrlh/Xuj3AYWB31qqt6/DcB1E/duLLHz9t91xPw+UZhh
jbOh9JVCOwcKNFeUU9Ey0ULqa55ciHf3rE7wAddbPv3yb1FZjMuCvvV3OZ55dZwtVatneb5NX4pE
fmY4Hs51zuBl03/SIvGJTvJMmp2xmihuk8MeEdL2Ah1bCfQ5lJFvctTNrzRaq6w4ixQ8QL/ZsjFG
RhbQQ9dwToHQ/bg7orYTvJ3Rzb9cgAROsjAMR02jKcVtdIQOqr/lZvsTgprI77eVJeKGlx0RCbtv
mfvkfhsp2vOv/JIJpwsCSf8or1LiqTjGENgp7WCgGjN3Z7rvn7PPQSd6j4wq3CsDuhCkX65Kclbp
TH+KP9FC9tY6oPzBlt+3N7aKW0s+Sd5uIZLrEnDa8XoWJmKoSqnCV0LC8dvEcFsBFS69t9ygmrbI
6VRE/pLFgLQ7IqzmXE74W/RVQVK1hZ1R5/nffs9xlYihVdxZ5OdXGnU6y16s8DI9fsWenK1w6pI9
iSoLFUoPRDWYwai/EuzxXvpX4LPXuqwGGoYF8CFb4RBgyXH0CqNU4WCQIuNVds/sluOQ97lTAf5I
msLfvIbENeQ+7wglQIXq1XZGrlyBPZOZ+TEZbycNspw/+Avom0LDXTxHeRDYwJwIQJL0ly82Lxgj
sM4tVl9e94LYURSwPHl+PUyLDENS4/oEfV10QFy81RWfOtTSDBFdVKQcC88fl3dPousOgORJ8TQG
hjvXv5fdhptkfbixfn2ZnXiPOpuu0nWINNWusTM720hDOvPnPfaFnrBTzEwYdJynX7/4Kr/Qzk2A
U2xS5ymuxjwNG2Y+P1B4tICx6/BLqtPAS/BmLcDgignfgk3OA28rnobjlb2dnlShyNbFU6Uz1BHP
d8UQ+OOMlik4Ur8h8mu7mPewxjAWud4+/gPqHeeb4dX3yCIpbWkC/6uYOAK81wkGe5pSTQPu9QV7
6j1HvFLPaUSuJSCauMzkdZSCztFcePl+VhNgrmL+MadJiqLl/hKLJHBHOkyFB4YDZQ6OGjnFWoWH
yy5phM9PCHlyK77zaS77DMnc25QH9VLrRd3KR4DHLlANb1kG72X4bmnzXhaaEWT1EifiqVsz+t6Q
TEHtIJaXVQrdpQg94Ndmn9SdTrhYlIv7kAh0CHuj+OdVcx97b+xqwlWZ2opzBWK+5ycoCwG0AsMl
11iKVpaAWgtph+l9EQUDRcMqh7n3Oci2vPwQIAX0flS3e3hg3XJesykDOjSJMVJG1fbYFcSEWMWY
iTrSoEGXhhuX6NJBLKQw2us8pdgYI9Ai0/8cSOJ2o90Alt3xbAMEoPjlx78MXmli+p139Luk5gl/
KTgoq3Fs2sfPjvNOlKUDG09cT5NW0oDXX4ZrGLCWnyyC0zGbkE89P4Ycc7jpzy/TpyvSGWmIZTtX
erENbJwqNbkU3bjKXTOA2hkZX+6rm8aiw/m/lvhPIPQthWPohKHZeq7qKOKd6y8ht7kLKsvZdrss
K+8rOrffH/MbfLK7YRaBxNdOfoKUid39ZYV9JPth9YYP5A/CuUh9O0sotrAPXFRwI3x6nbO5NpIH
DxBwh9ieynS+LWbFUeQU7qnibIsNIrrR7VYYH5r8kKtRr2b6bttyIwNIxEOqI0BuWsVTiNd3SvQn
mLRQO5Qd2pNHoDG9x/ocyfnLZd8InSjjUEwfAlGKkFk8ruYIBw3WTGt+1jtZnHWrjHiYN2uvh2Jt
eIXqv0oU10VvVinz+jwS+CB6cOGdC44eCTMR5nWm/6GX8S32fsvETHH3QpnnDDGlSuI4xqAS7H4D
beL2MKHjoXcVKtBZmz6J8xRvhqNKpouGNf5a5Lmx/juinzHtaUNLFgslWBhId2toDEUAfSHG/QVP
ytaJ7rl0JT9U3nMMdx8E0tVTtatcvsIypv0UgQGYKC3gWN2qQ2IRCzLRfrPpM1juB4Q+Vpp0LLfP
HEcZX1rbYdlxYMvTVj0xFCmezyAJHc3snXF4mqsFmi3O1NHoBqmZwYuevBrhh/pTzV1dXaQScs3w
199iBuvXUJvhysmA1SvlwErzVOgJjbCyZV2REirxQItGER7pB56NgVbE+uGdbSDF6KfjFF3JRd/E
H9mk60//OOw6Dj9vqEyemLZBg3Eun8FOGTYZE94P0FHaOPcDJoROHiUKVpWnbKQGwYCtU7vLjcYX
XRMTL7g8FSOy6hr8qYfCFX/Vg78KbfTGvAfH4heouLnDgR/k+p3pDaDc87VQrKiWXa1Ui859AXbf
nEY81iymZY76Mr5sXLsrn8QI75xoy3OpoQrEOyraUn0zhYee7wGt6YEZzTzMNRmvSO5P6jJSWp8O
Ibs6ueXs65mCVqwIc5BazzRoOdvSR+ulWRjHBaMH8fCRgs3O7OJ4/wDrfzCRbCVRWuNNaQciY8vh
Glb3WsJ7KloNIa7PiglhGCGCqDc4ZiR5C3N/6YL2EE2nT+vjrnn1mW8JLCXb9OYcPm088BlW6LOF
a/iQRuJKsNVIakLTaYYeSa822owmJ5ywXk9Ooxz/dFxCw9CVscF+IEQ2e8T71rgCwTjZ2UFrBC8a
gmdusgIU3hhfXT2/VBsXIKxts4JAnFikiJnicSiUfbPUwSkzhqgJ4bPMZcYQPFxkqHO9pkFue8Tb
JQBbJ3ijnd2m8HkVrfwiYoRyz41JrW+Z1qabCITQDVV1DhfMnUPeBGsART1V9Ox2GUHeLTakH06R
qhXWSY0pk5JFP29Xw4Y0TbOwa4DTm51YoJGc2Nj+d7qmPNVkfdvyzwe0am2OoMZjkEgZcZpfcNm1
cSfmxo9HK0FVAZd1ucyZzVe/99h8rBN2uUiHxh/mzm2NTFnVb1V0tlt3y2QSrfLjiHSrAPDzlcYd
6A+t7rBaFT/UCfXLchKB5m//zh+WxS9IewE/g5xSy3mryyUVU9UAHgxzj8LzFYTfWSnj0+hGJvnh
1Yh9mHH69VO5HNGJ61aFq1pmYq5hTGkFfKs90wnKArF7vfLs8unLhQfULUuU2P2o+q+lM9qeJ9X1
JrzZ4VJ11Peeeq/+p0q/hEz3soOCN8BJRysSkfeiKk7tCZvosDZsqpYLy12EIjfUOLx59sBVa+VC
EGz8Ah/WVcK6HGvE0+qSSWqFLoy+el39IDorX6VnHXrCPWhEIZWiZH9qmqzgFNqeofXk2oPFKYD/
nqUmTza6QanfGtugLRLNYezCiNqKs+zznKqx3VYU7q3pV5DdiouAO56nCzhDLuxjWI+PZhmD9bJk
HS79J2j8znOytoOpv3yaJavcWVZ+NW8mvjz4lNHayEDz6E9Ps6WDnneNf0XUk9w65DHF8bZMn/5X
JbXVkjBuz5hhOcnb/qvFru0FkRerb8wQRt7wrxFD6Tb8pyeVr0nLOasJcUaemhZLuf0XBeKK87N6
iJuf5Haxp/SAwWgWdPUMsz4NSmsi3RMGnNq6tIvuGACSgrPZwvpXq0FdNW/AsuBtNLE7iVaZxpOf
VFtapaeTa5yUDZHBFAlC0r9ns7iBs9tDhHzwIS8H1FafVfO2BuzxfePJo0RjzcWOzQtMWjrPH/7i
iagc7bUsw50eFV2Wnm/YqiqoMci1frTF0zq1fvIeKmWBSjAeVbk5/ntAkpAp6J+lB7sQoV/z87/n
YxU9tcnIJiDyAVyhh+fMBSCOb8CGAfyhaqAmSqBZlEtHOMDeS/EtjqZpULKDTtVowyULECWAc6Cu
aBQcEzneemXYQakbhKPyGDG1T/sRs3zD6dYXO92BQGxpQqsFYvMC7n/PDJpGA9H+b7+lD7Qkky7h
p7Y73jMb5mc/9IWPaI/gF+pg2R4BlfN5rApgKza0qJdie6W23HQq7RztNIwmpHMl/NODyrFy/BFg
S6xSJK4FMCHrn33vb0SzyimFN9TFvAaOXsc6VIHlU8M5IgQmk3DTTZCq+LTUcvJyCBVlAMXueqkM
nmROs1iYYeYBoD3AgzMYhymbAL3rq0e04hbA8CerBvPY71u4a1k3kmgW9+I70vMZ+N3TeiSMf11L
XBzwwabyJYMi621y/fBiQ+tiAcSFYVBm91R1uCH52zlKdAI7TSzbtBcrrwqXpl9MBq5ICAciK1wK
lMe5jYrzkeSeLXjh1WBftTRtRtgYqDlM1Up1f8ZMXL5rwoFJGLy6VeTN10IwsTB5HIcTaSQ+DppN
E1NtUI1DyASuImXyuYioPKRkixCUuzk7jlmiKRwEHfAFI94Vh7NE79VZ/AgdnAPeZV7zG38Esuwa
6EZtYH0ey7FPiAQPiBI4JTb6qyIXxmU+i350kS5FiJkMsMHufj2eLT5sWaMRmHfxBxm0yVNvzpht
gpVXNlg7PsSkTPSaLUmg7oGJz27xCpjf98pvn6b+FeomvoDIMIS5o8sizCxm4c28m+SOrs7hOuPj
p8TQULDVYQZO1e+cRwfiahvmMYzOAdy0W3nfj3s+8HWxbfrZ33G5RqK5J8d/i/opC/1UFS7A0LWQ
GwjkIo/wLNjGA4O/cgA0X0o3uJGBK07yhS7Gqdf9ptY+lXeetykw8nxOPEA2MyDVSut++7z63i+3
ukP0Y6q/y0jro6GFSe9FclkAWmOoX0Z8ELwEXpleDH8/IR1FDHiYgMwyAPVACwgnENUBfc8yZi4C
1EJu8vaSTwsuTQ9Yu3Xyw8+QcW7Wiy+VGrwnvXALASbtXiyb0+/GkH+oCSWJ2d8O0IPcIYFUj1vT
eMErqQOIHa/UlLi+ndBY08AL5+gEojkNTlKqUX6wz/LQgFbpgL9B0Knyavjyn/BMB89/PO/XdlbU
EVI8Y34/3/VejVASHqcyTJXPC9yod64uLNEnFm0QM+3CY4msraSHjjy5GOO4Ls2o1mWZifVoykcN
VsIn3x7VSU5NHypw+lV1xML5oRAckJD1UosvCsQ1lKPtY8oa3wvcJWTfyQIpxXk1icD0dbGjuZb3
dlNHehrF0o+ApTSUI70v3Owut3VOpLExVhePyqwP/RrEeLBTouyx4cleo4oBCMFpLbmr/yvDV9FI
JZ3Vwk0FAm9l7fALtVQmG+PLNmC0V9GPf9uCmGztg10D3sOOzoagymb3olTVsSSF3+kf/BwnOYuf
eUYQabxiDKEepMYH+F3wkmgo49jk69/vv4cMS62icmFuPrWkBupOnk6kn0tezsTdGmZIIXFv5L0n
FXcKwyA354W4KMISYyQuO7Xh1trUmkeZJkcThqwnuQOjVAQurr1P97fL6k1iQ02LsU55PGZmS8GY
cAOga8KHBKuan4a45MqHUty1fkrx7M3I/iqzN92/WXGYXPmCXJRIzuY7K5E9UAL/251GXE3pUoBo
CSwr097mV4JWIJloRqBtN+5w22q2D+HXVrNSsKXq4xF7HpUgqlCiDvoCUf5OT9NyRLbM+SEBM5xH
3m/diTPkN0HcCKRJxxjDe9SNbLec9FhAdsIPpBpa7GNXahuzJGIhERVDioZsT3kBsBeiBIxDyJTr
5VKxrNJbeB70nMjwR6O/7Lgw9FdDHMX7eMEQiKdCRWd3GpzoJhN1gDntKymBhkfJCwiQvlZFDGGx
q2X2Tvfjne/4G9LCLj2/BtS7NaOLWSYjjEgPaFgKh8C3Kdn3r8uruBuHW2U+ZAdXEHrOSolwO8Q1
bKML91mHsSgik2kHM89AtwhKXh/XIkpjTHR/jD+ZS6K+l4Xl5M3yvwCNPB+CvUgOA0lYUk7p6tcn
EFqaQleJNrL1Sk/1bb7Ea1sdoV2Z/66QQeYzHL0RVdEmRoO1CBv6jAo+Ij+FBfBpZJlJqr4grIRJ
S37vyW9dH4W6BOshZXwTXeSH8SK0j3isI55LUeqnQtuemoW0qX7o4wObsMzGZa5LmB4joOG0mTmw
Z+iXbzUPQ4FcKOqDlqNaGA5o2GyOmW2ldot7XQ2V4D8spClUDfTjYWQzG9C+w7oikQLnXK7HuCm0
S3vV+9N7Wc/K+QQsgGFA8H70haNR45+rqd9s9gzRMufCnIJPiO++jekDPbZJuRmvuXqsUa8TlnAR
grpFLewsQ7csZ5IZjCfPOzjQM8X3gIqsTY9XkZWx3uqwDzZOMZlNL/EUCgMUrsh132ScIlt54yhK
kPLStN1tEydsetI+9jPe+mvPNyYuIuwYehBmpqGPoPQH6YKpKEfPVYW8KCHdqkm673w8INKRFKdg
3oXqp5ulHW4FbCQlL93ejT47o1RMXrof7B5O1pjJk5HE7xEBxy2UJXx3Ovw7Vbq3RAW5GGQdc/7Y
VBQAZc9wa1LjpjMk3V9PZYY6aprWIlN9vnWAW+F7vx9SKm7d7PzzUwgrqg1FzFwt4VL3KEHL6NsX
M9VMoY52K6xQuHh7wq9YaV3fpNRcSzXSDXwpPPwYSvbQqdBopI6IdMX7UqfP3/W3VyV1FQY1cpki
K3EaNYG8eq9CpACVOcEYiVx/am+efhQyvW3qzfs6S4VpTa63Vo7Jb6BSldhnzGrsWFD7jp23909A
W5VCdA/pLFd5IijoNTBaOTho5HX5KMHdo1iO6sjpkvSbYHz9tBD2JQXfo93IL/cnjGR6r1Qb60UX
DWXpg81dF+ez84KaIS6OFUrjgME5t6+M8M2dPN1CYBdfaHyWIS0e5Yeb36WAZLGRqhhMrTYBtHTp
ZMssHBDwX4fHi8tzB9ofUm1U764Oj0zurdVQxtpI6cmzs5AxUdzFfsVlO3fUEjWZt3yacOi2pht+
Ry8B9+SrY9tk1l/JddiLEk1fT6y1eI/i205kfvVOMbxJFS7bZbZEccLVRiZq8I7HSdX5iersHmpv
hDGodY117UG+MoVr9JZ2XEQYABIAOKnwI7fGGTgnOHc4hJGRXn0yoxPtRh62OGyImq++plzMNq0t
DMwwM5ZOAKJhTtmhKDtI33SURsrJZcsger1IiE9RSxbVuMWgZG/yHh+XICcWPhwOgnKZhHHG6/Bm
9LkW0zHpOqcqYFq43b7sp+0j8oyLe8Zq6SWhyLb1E+CF0EXzD2TIzWFijRFDEK2SGWUHg2LBxeDd
RBeIUZbdmUot0h3VVB9NXeKAyK/2Viwlm8pFPceM5vFuMoleUSTfxGzRsRTRrCiSDa1XI/hlhHT8
IRD+cdyVwBhHbvIqdPCBoa/qZQJAtjolgBUG0tkjYT0QJBJqESGS1cvvJSorLMDZTV99NMGP6K+X
Qd0qxkLlHDDv4LttgYKJXHyGBl3cvtmuwcLLkqcg31yRnlzwnl3HrlTV8wj8GgRHXE7AQYym/uR8
kOjJe0NBKc6pfomwff+ThUSoI981Gh6oloiVy+rtrGRS+dWoiPWsbHk5Oa5mdzjHKRzsub0sX+73
yg+VXIg+lIobiXFxUWgNbcCo/2UhfXAWYvEd95k4dn2vIiZD59eunkitj1ftAOF7b5xZj7vsZQ5M
ZoYH/vr9dbWCsmtqPM5OYceE4sMSq2QiQ12Juckdtd7FvcFl7+O7cz0tTtA+zzezm83EQDa/JZBz
mSPO2JniEhPnRmiexprrG4wNjIF8qzTeptn80PF/F688/nY7MeNAr33o/WI+OAm77xzRqXwzJiwu
vVHfByJQwQlsDQM8thR6Ep/Iz39RWFeitaFkqFW91KnSz9clab7s9x/gE3vxScUNHwToYkDCL+Ce
FD6xPIAJRo9K74OufhdX5G39uaA50YzIqiYR2WKzZZwHEbk9SMfUR1FlaEnQba2qChgDrSItOX+P
pPXekiumHl/iynYDmzWN/IvlajioNYo5tEA5XaaFDmzJwqM+d7fJ2Se0Kfszu0Ef5WD4FCkWP+Is
CdaWZrw+FcHVzW7Yz/1u1AKZTJWhIlzcFHF9HjAimgAEUZ5Duhf/CFGOIY/V8XHbWGdUbP6it8Em
Sh513BOVuLvZzJHh/bpVBAjmu5LGaZu1t1bOUKVnXFIN3KLd3eqvsGL2A9qzMXgSHKB2YHhf+ZuV
CTTXWCzFTRwnLAxWwyHx1ONEF7hg7d+ryxE5e8vBKPgCAZJPGb/FzJbo1MRBBzPSPPEsMEQxj69c
KPFabnwTmYuLQhwlc8gqGC2v1An6BJomvCuFZ1RdRzag/x7KK7Uefjxc1cw45X2Og4H75hsytKN6
2WbgaGeTmyrm4yLWXwlioFVyPGLjFTPizk4KZEv20nTHqBishWidlH+HIDhxFIXHua67hfMICsP3
8n8g+xDTiOEfKvVr9zpjnaglfm/liSFjJAXU7WRA9v8csw9Nej9Pjj9OZ9VhGClqgf9FI+4VLjdc
4yy90VjGrFKdAxhRjTJjdidQaMLGsRu/BULgWww9K5vHOFxH7jRuxQ1KkxCkzNoNrTUGH2K591DE
0e/hJafLzQw+8WvI2TMtOH7e8xE9xMulHXrYyKZRCQHZ1REp4fBCg7XU2WlcHogBrPUc40ioNPD5
SpJ2outjREkte5gn9VtibJWwSR1ibU1pJhPoWJWMacySDl6K8UAiQIwppAE6MvwtbOmn4rPHmAso
Rjv+99M1GPmNYI7CrXyMrw/5oncQCBn7KUAqz4eCJu7erhh1eZJm+rPUdR58wOeWJe6/TFyOR0Ni
FGE8T3SkUdNtOr228JnwiDybBXumyKWUDisdro+wcTJYPXTHueLrBVbflY8Ob3G+QhG5EQ5Lw5PO
J+rcNGDN1arXX+lbAYHiIrMTJ0AUiFhjbdYCAP2/JWGUugD6aqgMb3dYKSws81OBFuEyH9wG5xiq
BUisfRpaIpIV2eZz7pkrtJkj24ejHibqGDDAKfPY6Y/fsM88gtVfPgxV/P2ncjmNogC0R56vTiqV
mJoQpSi+n7XF5Pw/ZBQfKagiU0fnBqWj/qDNYUyqB5myunDvyINsTXIkSP3d5J/XseEI0y9Rvdsu
ROyNC5yDhvHzhYGyyBEgtF2smlv1vqo/qgMVSM2wnt3/hSEcubxr667/RGDx1/4abPMxcf5SFUaF
V9pW9ZRyWM+2m28RAv7UzLdvCGAl1jcM7c5WQdOAnUiJVcsDSHE9pdcm9XMlhW1+r7R7y41n4hdE
geC7EQxvykhtkyhTALPwtBWBGwQZz8t+snAmZ8ANPIsDIOtF2iF1UF6uvVeqgMdm/4z+HA3sH28a
U+GE4eEVgZ8PrF+7nF0Zz39HHcYllM7RKY/DhNnUrg3Jpn80vxhN1gdk/da4ecxLpTWMntqa8Iui
5kLM1bessFWIUXMB6seIo9bFL+meH1vuLsDnv1oduKGO/WBdvVc9Qqq3ZKRh21Ww0SYoWqN+E5vM
b3Hu3sXSpEwObcgVgaUv5dSEeGU9Y+OvhWP7B8sQSShc21oyk4iq90tv5Fa2yJmYlmf7uaytFw3s
pSjGrQ7/fKVt0qLyRUuzjWnWMouKg7bXARot3uZTGb4K8GDCSv2D9BWkcwcMfEIs5l+PS5gVSRle
MJNS+q1mCNMe50JRrO3wojaSQhhhNYf2CV2ovFC/6WiNtul0WdaZ50FW9xcYMP/DJGfZdM8jr0SA
qM0MGARcmLuvMYtIuMblp3CsR5IlvLRHQuzibL72Hznm/0z89XxEzQH7IlElb+7jPKNR/jpMvJQg
xxfAyYQwUxs5ZlV+ntL/FAqmIIf9Rzq/WC69gr7UoNmIzfEqHyvDgmBTLIT1sd3EBowlGiHjbDNR
/dT1RwXWb5vh5kZFxZgNZjTAmHXmYJTZa0mebBBJ2RJsw/LePYE9nofEiFklv3SUWVu+kkeW6xIm
F+NyIlEwr5/b16U7tMsE8f8GdGJ99HSn6mgKB9L/fv7O3oDsLWkG1gWDA18KN8gQj+/LgJHNahcA
xoSO3FpjINzFc0YQrXHIX3E/ma1ZNmXWUTo4aDAI5hj2RmM9oVtYGixcyCxf+Nu7NcxPMPWwKnCA
Dc2nzkwqI9e26arqlpGQELOqTRo3t6d2Me7hrhSxelhAhceDAe2OBQ/EVjTojBQ5zcI03hzzAkaG
o30C+4mOPFPQGJwDrUF2IO2PM+XWxY6wmNpgdl9bpfgcSyUH0vlybzv8ONhNTYT77h7gyIFPSj0S
g2u0C6LXU+JpCzv/594DOMGci/s0WYj5ha721ZUzPoePqIctCPbWAb5UeuOWll/sCyM17Qsb1h7m
jGMkHpeTYtAbBkt0kevXvmahnIQ2g+eKjdn2AWFuWF10xINozNF+dhAC2cTmHy7sWkawwB73p2T5
zLrcIeFVvxWWw5SmCkVaIiircAGwLXFxBQfgckYEiLgpMSQDtKCHYFAwnwxqZJs1iEpAHBD0R488
N4eWStfebnFgS8GSKgKpr19v4DM5iaqKCPpeIeLsmdCkzCF88Lymuxtg35opna9iHdzAM2afly1R
TP2Fq9lM2xNW5mh35CSsAB5wL/X1kAVBngfq4g571imuDLbRKjEW1d6ofErRlpvxIdZQyyh1jpga
zz2l6LJWVEPoyzd+VwbgG+anwtyyolnZUu1JdZAwCQwxchBFWizl9tuOSzE1OrPu8pjka+UwiyFY
TybEUIJp52/1NjALxyFyErGq7qofrYaHGkjGOi6syOhQ0tU4aLkLi6U4BfIPnvAG7gdTaOniTWfa
tFn6A7knujXrt4+ExcnLJ+B/metn29AAXdOL/OO7jXT5sgsEJwCNmevJNVvzgURk7ng82Yfj/xTj
sSfsT2C1F5CZrsLBcxSfhTdbLekZvobCvmuEGXVRd+wGo2v2Cra52Ln7XGaDH3X8MXRfy+zdgalU
9wE/zQWHKLmI1XpI6lkRn5A3VuIF/9EE6Ha3+QM6YJGomnLoDM/QOKCYw4rZrSvP6cx0eIuZHe7q
zOHNwB0wCOmoxmc2+dG/1pC4rtEyNWwhZgrp/y7Ohg3Wfl1z6qDpdb4e2B/Y1S2b+h9GyuQtk+9A
PjGV3c2XojVtOB1XnINg5BJCPqTCBJ6rWtzlLwG3QenNeBqVq0VwKcVgcFk0cLWMS7mUMIafYvd2
MqPHhzlYhU0DNGA9QSIyrhc7MnQQPmom1vdX/6azC8A3ccxo+PQZ/1frIkAL90xcZ2KloTPIoSao
So5vd/OLiKtnY/oUFOQfawkH5U7Mvv+kzSwpYtldV5loU7jOy5ApBrXzayD3tqNbTHJCS53Xp835
dKn1t8YnMDzX60DiDkzJjRZlZMcksqEv4XRMcae4Z/p/vFuEW+2+sxhn1iIPtXcq+BMRfqs7wG8M
NaAmSAKi09Pqvg0UBHhqHs0848s0JR94cyhHW2qcHQ3JWxo4z0j+m4Zwx+t/ic97bzCt76LxW8FZ
yYw8N8iPxeBuoeU+HIfnWWtnM4fW3zKsnTdRbEA/RiUoLmlF3vWCe9Da4wfSspmPmLJOzA9o6bc/
JvUOdY66HG9Mrj4Ffu9uyjpsZRU59gUbZbuNSbzlRjZUn+XH/5tpvIn1+FCEgXhliblu16xM3FKC
a/wEWt8/Z2wNvMcuXXIKScrAbT7AP8uUe/SzyR8vBq4hTJuhxM/9ZKvckot6KqxU6pbIqgWo7Bz9
WUAtYYrUZHdNqPOnHYmt+AgTKtlZo/4xCKiprWgKpj/dU4bpMfu5m1mkjjczQvmdxzjeux/Op4v9
wSKQDCEaK5+6yNZAiE1cAKvZ+K9CYphz3WWJq/bIxXPw7z14paIW4TAPGQ/Z6yljPTxQ4BourFWR
nhxwE4LDOn3iuHlRBPlv8/YzGtEjPl3uQtml/VqEpioIWOgQCUCqoEmR24XLQYRtRrwqYAHVqArO
vUge9u38ugMWSoSX2jgUsbkHJicwAqxIB3clPrQCSJyZ9iyLcfUvdpMXGt/8zJsxXv/zBrjDXgtg
5jdRrlLW2gReNMxtRgI7Xq5XhbDWt/XAE6X4aItSyD+2cLEz5vJ+yqa89LIwOQyh+jy4o5iU1uSr
pqeIWFWSb45RzvrX5W5kMXJWGZwcArhRRJSpTvbeXzIUi6027VwGKjDNlI6gdO7fwUWoVVPxA7eB
NknrIRpdkc8BmopRhtaeWKg+rwxHtnKHFyDzPmThj+h7yPNHoBs2anqiUL7o42SfzOKQIq3yEau5
2Dm5dDRn2Z7Gjt4yQNye9amiS9Q6ulRN0ImCAosQ+P9QTZWEmmy88JhuOkfIHpIWKEnqx/IEXixP
D3fGvDeFJNm9PYdZ/8yQBvrn8StqLEEn7ap0pyrSHgMM1XdtF5eP1BHs3tWH/zhFmfPEyAO3rJMp
eM7QDtfPODgAVTLNl9pL2h93tuATV9vNu376EtjXlBMSYQOZExaOFO+1VKSZv2QlMtbbolH8iQK2
NL3EDGhBEOAjQ2F0WSsvGku49ywBBLv2EApm0ihNbFEhA+v/igoxNNj4DVRdzOq2zkIZK8FsJWmt
uT7YIfKJ+gdeURHDijN7bXBX7Vza6L3gtOBJkj+bU26T8Kw3KaVkZP1gmhpRxKkWdt27eCz2py8y
O5cl8ShV/0gHLW8gXatQ/gk3WNF6qCy/uF5LgifE9i/82Khn3aH3XyFwDLu0jNSe360yW1L9wBJo
b4cHebxpckuKHtvZ4hV3oS9+6jw3JikV0m34HUUaRncyy8w2oV0rx85VRmtI3voUSDrjwriFW9M8
qNfLRSJVo7vrTa3PgmmVeQD2TFVOrDNhesVkAZ1Ve3igWABtIDVFQGgnvAUKrP01HjBlC9JeLhwG
v1ZgUiBNXz4/xi9JFY3pMOdQTOn+Y3m7YB4ryPHxExTnHDDe80UjG8vD8EV3t5HQyFqnEIAX8Oi5
LgqhBCMaTA3Xx4x+8GB6vSZ5HDpAiT1/L9n+oIxo+my7s7wO8NFOHqxCKwi4bwK+usvLJUAH0UUR
KP2Ry28+xHBPeDpNHcGcBZlVfbDZe8U9c1pybPFdAU9dAIolfgcKucQkO8yyvlUiTWDWi5QFwXms
bdcuytFk/Gqu8q8xiObTBEhMqUZYs/EgL6jwGXLeozsNJJmcWdWgLt8Ec5u+P4DF7kM7mkilV0VA
qArlkWU//h9HyHGViuMxVhaMdRXQI3vHT5JfC/LHwddzYh0fVH21VodMcensTYUtoawurfEDiuaT
w/EZSVabTAUA4qW/zd3Xl3k4HYNaulWL8u8rWaRcY5yq/zKmso46+UjXnceHnoqs5IKAUdfyaMDz
sGwJ5tZOGoCxgpU+tt+t2UU1ZdZABNkj1k+RciXmzM2cDgPDBoPvcfowM3WP9TWs33PaqEjfVRCI
mvtXl8k+/iOHQW5RIvezm/cA0msgv9ps2meyDfRsWfTVSO/4u7nTQA+B6h7e8PafwfV5Vso/s2DT
k1pAdo25BzRrNQObYQnJLslC4/uEqxcnlicTJ/fLamE/AVs5MU/p90MNxaDnjvbNCjTWGQl4aauV
M+a8TLUPvu3EnmBerZQKdNOW1+QtTjAa3yMlCVY8OULf0XaRIcnJiAS2idoAnYHIsUEgdFGMmicr
hUofHzurdG1OZJx/d02bzvRbX1DsIXmcLlJTgMe0OwUpJwTvGIpX9LTNs8xg9Y/Sn1tVDwK/jiqn
rZ+RMq1Y+11/0xV3ooGNzCLo5P9kLk1VEknoKh6HOZg5PU0BG2POrtkeDjqvY0nxsQ9R9OOL1FaR
zRNUkkBdeiLF5TrgJCzbmgvI6uo0mZX05RsFBagNdVDIiPY5sl+8yKG07KWXkjAg1Us+AJUfM85U
KvaVjRIXPKEeLH0cwBNTyglvkAwNQFbsThtW5pAbXHGVSaW5OaAg2aNSMPH6VlS2c7QqZWLLCcu3
aUav+moo49Mg74T9sUsNAyog7M07n/rP8VsoGTfAcQtEy2gXXgdoeTb4lw4CZ5CeRb8h4XScvVfZ
PAoXpT642j/an+r40EGS6jZdEoCenKX31om6ZKedHQBc2S9ANI5PYDG3KJS6NDcdJQW8L5xEtTW+
E9UmtjsI3kRlv6Ysgxx/m5ktbfIQZ0Br/B+nJLHWIJ7i8aKMa0mGtFzqGf5HhzaGcbL8/DlUVtgy
s6JrHNHsG+yLwwkxnfZhIU/zJXMck05sVrghVr6QnJgg+pdh00PfvzdBTB26ywrvCC/sZrSE2eQ/
TALAA4PBNBCCSJ3GqC7uqIw9QF+l7fs6+sxNU6Te51XAoFlvfgPYKnwKFLavSX8S+TVLH4WjDRXq
KcCGRvPl/zy0jKuukDwoPVoekQ/CrHtd1GzeLQaWRdQ8SvJA0QzS9+Q3NSyCMZutlnL0LOEwR4hO
l1j+gi3EOEENYzAk+4nllJ4fCChdY5kKWQN87M9jEoqm0fgSRTjPyDbEqQEbPMR97xoF0bpCBGLI
wh6nSIpqlqxr6Wk4m6wbp9/xkR6SP/vdWH7ydc6Z3eBV+5g989F1d2/m26a8o7S8hA7xTGJDhPIa
j/b/ZyOKI+PWu36k6sTrWRz4qEJovSdSedbM7d/u4aK5cvwVnYhRWq2zb5iLcGBKl++EQSni0mRO
RfeB6TTY04vf22Vd8Cu1qJ9l/PtzSevvgYgpufe/kYApnSSjLSZwXVDEGZW2aZ16FAxtjEyX2zyX
w906TqD2ohU8TKRPtirZGF54S0nJFq0lBSAbhZFIz9lExpj05/aneQqqakpIZhZZ/qBk9kCgEljB
diWLoaxuVA0aEt6X0xU/x+v9M634mAf4f7wGTtCY2roF8ANvTg+kQjAffAUjEYQT1ggrGEgg/0Ca
xZJEP6+VN9J3FZEIScbuyDU9iRB1ND0k+oqag0pRz25ORqZQV4KsQUXbFKnbQ0VuzDTf5UQYd1VZ
GJbr3Js5b8z026LB1cWeFbVUlDFb8kP7AWKNBIgo1FDXFpGNByy4UpEmScoJiUgPg0QwtYcBPgOg
CyLwFY+ZJl8qOv1ZCDXHtrvPtNHCOETHtCeRnLQpsr57bS82nF2sbcVdH0YWUZ5taB0IYUA7bWF5
/Hwe00lagR/1qpGRSHJNi/t1cD75Zn7TfYMAirSuyJ+12zujoGaDF1EWRwgG4OZpI4uzntJLDoSU
7+HUR90J6fOKUCTgBY6OpMJaqrCbWaMv+6BYPL2DNYk+VPc1buLuZAVFt8YNwtYcpTGseuemqsXu
HulXdmAI1QQVF8fdGYrK6fjIgIEt3dUvHFbJ7OHWXtRq3H3tu6Q0VSpSE3C1e4NCh1DXdqMyuOmX
fBParX0qoTMC9iORLj25ucGVD+5zzzQ8UBXLiFD6puPVRi/HcZ4T0MKxOtcNfFX8xQRlZTk9vIzL
tzRHjBlxw+ykwx+1ws/ifUi92wgCKiRxx2PxkC61UqnTPMgeHFWqtxNURCiZ0uiCPvczl5EKv23q
2FAkvCa9SV+ibKDFhYXYtMODZxjU+xE64bZEoSW1cY+4Ngyr2iKw3DwdDX3U7q/yNOAlNTryxTb4
Rei4n52POeSgSiPJHwcEXbrP9vn46tyYnwU05su6BE+cm55tJm3WfH5EN1U1s0JAnDvh6UaXS3xU
DEWUfWUVkmdtmscZ/0iAktMPZWb4jxrrghxlMRpORYpGsugC00MiTJ8Kk4WxC/shzuvjdTZD9M5j
aLGN91UhJMc2kF2cEVtQGoFjjJkBAtwcYgl1X9cxwXBo5/yVpQ3xfxJdvQlNIbxN+GGHQLa3B+1H
/yM2KxbcbpO++7IpQTKnsOSr9N+mw7OJG2JIPAH37x0jeLhlW7pdQN6HKs9O1XHvLwM+RAG4lYNB
7SWNgU9ZoM+GOz/RAc9CiJL5XFAGpB1yE4eGzvXHHnkCmwNDnxljwtEOTZVTAHgr037p90HPkn83
c2aLTwJ6g/Qg3QkgrV0BEbgFgeNmmFmpGw0nUBElTBgGb0glJXAI2imy4tdjyuDsmysTHnIXqlaS
SXIjI+d6f4QxzwyYsz6/yV9JEvvu7UlJDYxA+ITi4iz1QHwv0YHvrLrpkj5yTVCbgU54ySK9LPla
NnjBgoBajZHWLP8FY4+AoLSf3NZHx7ZaLXBUhT0GfmX1ZVUSW6jmDbBr5jXrzE5uJ/WLs5F8RTrQ
dtjbriVlH7mfuqN7AqESswpDWB3XeKI4Qqn1GB6S15nPwvGCPfb2H7mzF9N4wYwtTScWsctRUj71
8i4lvj35oYOCtSIvGBvXQ/Q7SEPfT8MudanBcYh/hkUWU7yQ2Z43El8h+Ugv0uQ4SAfjfbpaUC/u
bGEvbh1lmKwiaqLAZn4TshvwvpXBpF0h76ynUWPrf/zs7M7N8d3Qf60KCUJ13D19svNrLloSL1v1
0IJbfgfbeVdrZ5ODWzJBHWELvJjWP0x2EgorG6H1UVcARkpOAyapevDwQgCH90rk6WDOVTHbuLYq
38jlaUvjXtt21Hepzu6TbuSZ7yXe/M6WLcYJMgUXfmN64GPJUyn/I7GhPY3iGSq+HeX5nf05HJIJ
enb6yQev7ut2DcHkR7U2Q8KntbNaNbJej98jeGri6yDeoQkMdDtL9oGWfhsVNOivGtSD5lhENkgu
FV9ndTAw2i9keD/O52LdgR/CVQqq24TsMCpjs1u3VPHf9Adl5oOkTugGmhh4ZE+APxKcduqo18ps
Hp/ztb20ry40gWTW+Ac4rs5v0Lb9fm5K+ERTd+qBQQEZ9Gzrfa7KoWdzgpQqRaWQOBRrlTjyk0OO
8bvgbwh6NiAvznNKc8eFPJLtauo1G6oRflR6rQjiiveLw1UHw8Z7dMddw7wp/yCSdgpnTECYWgsL
Mo7yXCjJX0qcnyX3ZtQ1DWUETYJw2ze14gr4cLbF46gcj1a8D+606keimq+pcINXoyoCJyInXQnu
hbkJN8izbbXyfRxDJIWnZgeFwKRA3ISPYCOQyC3IyBeyK5pk4u8al0brD477F3naUvD8mahuJ5ps
kLxojn0kUla42pbG+cFXqATsbulpGKvdL61qIn5H2sCQ2OwsOjGF+rDrFVi/NqSNWDB3g0Z9RkEL
A4jX889iqQT5k+Y1K7bBwr2gT6+bqbg/bbnH4Rnl8uqFhx9zpB1GF6WTOXn+LcWVvvVqgU+6r0kw
7XxNAfeNIFA+l2n/WpHg0XO4iHYI8zIcgdj5BvSiYJc1WHNHtiZAibUYjTZlnBQGTDT1/cfpPfaC
uUTiZlzaraXywuK1O6YoizV6j47chlg3sB6bNwwliIvgTGcj13gSITbUn11j408KVSed0xHOI+Zm
PwwiVLDUZeEEvIGZPmxO65V9OR1cVxJwNwEcn5oC7EjLVlOHJJLwyLChkfGrvy2ZGyU9N/BSF6j0
ZrCq5F6oPi2qV/yegmN6uD97UFD/phNLuWDDcnd0sT/N81uViUOEH5z9J3P7w6UcG3piR7RZgS8v
/2qfSZtFatqRqs7ajCxGP8Zh9XzfxHIxbwnoIBEz8vzpxy01v/OFreBI0/6DYeF/24VhAVIXvBv2
JcXSemcfZf/TrdpxAIKTagiBkMlqGKMhM/Krp5HpN3O1AF4DdQGO2OqneAr89B0gz/1m2W1pUl45
2pl7PBiNWX0Y1p4dVug0gbScoswSb4kpYzJ1CD0EjW4p7c6AzSBhAD26N3+ut+6oEGY/Lf2LsWbG
YAgUCyUq3r2zoY53kqHkjHb88RjJj8wO1M//yux12A9sh6N+qzoRipjCz/EshkpPbSkAnv21VPRl
oz0HtLx23DAXPQkTlE1+9m90HKmOQdAF/cdqRp6uvyPn59Coc8uP4mbC4Ykr1POequ/10kc9/WG7
Tl7+3EWMGc5G2MV6qr41+uhANN2dm5yW5VqGUPJGUOZULnGnjGOGjpWZKs2yzISL4oStBk7E/ASu
/+8bDhMoUzkcIeTHyBw05/LLVh79FAf9cwfJy/Dbqh6kL0CltG/hfR0PB8wVFXXfKY+oEPch0oV7
5X+a96s4ttmoqnsATbXXeDSUJVPYEVpbLugIMZ4Wj+Oe8vS561fVI8GTcsZQhJ6sa07uI0IDXAyg
T+5ti3B9TtrVhjQrUtf8/+iNA9DDzTJVHkXJqcjC80kipL5K4X+DFAMbUorqcgziNxtkUOUnX3p7
lZ7tT/ExnKFp1MI6U8tnulOf5xd8mLzd/lorm3g+neGVdjh4immZvh+XUfMJ0cfH54lY5pelRFuF
on/zOwcX1HOI5/Syr8siPlozgyQwLLULmZf6RZ5erQquhGZjlC5LdD31Ljg0MI3h1vektmXbl/ZA
RWVctWeGJEX1uUbYudjZw8x16+a13bKvjLVnf6+DRCjDv4teImF6NhI2K+5VTXSMsmyaCq++KtHc
SY9hPd0DSHN0DqG1db7M6QQTtHO7RprRKulRp7akn2yLfVaT+MualSWc50JXB/cw6TmM0qE6HIHq
9cwusArsTdZ3E2Bdg52mAW7TPVGg68IY+ijKhGIsgRs0qBGBEyhianxKE9nfzF6rkXKoCm7u2eCd
ChI7ePoRY2EGX+0o5ibDTKfn2x+Tq7GYxkOK6uzDZkZ6o68DYKf9fF9brX2xvtDPFzacPypeb2YK
eAEQGO2YSr70msa08wINyhD5aeiPwtXEONNp8UMd/TgQW5V0q/SYy9eiOqsFfVkfWAW1KDS2bsJ/
FInjrgtEP2EC+tSQ6lBqXJ9BW/RUuRbMl67xgtp9C695TqW0DwXgqQdyzLdzTmERf2mRGw+Cvz0T
a+7nj29hn2nT0Y3oGRJMEyctTg6EsBB/4P6oPIiT6mBajgSrwAwE2+FRJAirQTVw8EvUdpPJzQ6n
lZt90OPacERqW0CZHpP3Ok/03IRv0HAQ7U+U4J7K+4/M1jzLQXlq5pfeTe/YPiGWqX8UeIB2cmtx
mdv6rQyndUrCbGFF/zVQ3odcw17n7mQI4L82YKeExn8J/PBc51hFUvq9I3rwf6dMWUW/vBIh9iq6
3LyPnzjCVk6wV924ewCiE9ZaXtsw2IhlZlGB452zDoxrv/jpb8VuxBzY7YrcsMvSQZTsIq7aWni6
JKf7GShPh8FOnneHywAM1hjXX4Wp0RUkihCeqmpCwa8aX1uIDWS/VNy292+9FNmwbQREMlPOFgkD
m7B70Q6ATeZYUJldbJ0xo4uWWJtp1qsKiN8EKDBmacHfVXwXiADyKygBOmAJMmOgtAtYfp6vqBRX
r8n4dliBaS6H9L0sO1Jp5fO9tRXAxIYpkFYau3HZvus6GeHy5K3a4Lt++m6msKc1UWKYpFMXgD9q
ZxhJtQXNNKZFOd0rnBnNR86uetj/WQmEOCqZwftwah0dbE/RvJLZ8Tcbzbtx0WDQCzjh5De5G668
fkRFP5uCWNu2txGS2mFL9XB2xUpIphj1XijBFfGXPDhMT/UqO5MR2QnyZrsr4YQHRhj2TRlBB9BJ
h7TJr7phYRaPJs4B8O+NK7hYAilaKRke1D5oQN/L7ErnazvqiEszOx0fdi0cdYOZ26KoDaZuWB86
3KRLklhhYcGqnxDBuBcoMQDLJhoTx1cuJnoRvHsdj7SVelsG3eNx+YZlDgBAsRl1NsgfMZkgBt02
ewDZDfn4+wJHgKXeQqDhgjJQZH3qrfRaFZvzwJvptvnYsZ5yrQ37hV1hTCkNm47iOl/tu0OiGis1
frx0Vp+IzXHZtopt+QTDCjysjznSSO+tty1KfnNTalKkCh3jf6br/0NWq1JAX/MCIUjzr2Lcx6jL
iJRHyThKdf1aQt3gHzH82kluWjvhJi2I4OdklLfLKbcTpFcTn9jM6kmyvdSTgJZ2TmK3HG7UdU7u
2e69dnx5lr9iifCmES3MsqtldFWJy1jy8tTzYDY7g59xB+mS3112BiYGfNaAycmMaSdquhiIdhVS
zZnH651aF+vtT8W02dN0MBdOhdx7Yz68K0Pw+4Fkb3/V4Mn1TRpif5K6M+7qyPFcMPxCve105gsn
TTtx0YapoP+ZV2HeUA4h6nwMuR1f2vhFALqHuZfH2bd/smm4blAfEHq0EZiH1IQvUHxj7Ri2G90l
/BMPdB4DaSkcBxyfutQNs7ilB5kc92tbBNUPCTfVukzUU+vTndtvVmLJ0PX+OMZRFAbJMC2XS9Ax
aF7rmi2MpzXqZBU7GQYhtxUNqqsKQyQciFrEHkhtibARUI953I5pgEpUbbedFqhLpylYeOcGUyyl
3KGxe/DiP4xfJbMhc+EFzVxrB+jnRkTM4Ed5RE2n4UmOPV0XopCSnI+xw87+sifJAg7MVN3nu2Hh
AXs89s28u+x2irLiWEIu/N3Wt2mPm860LLAa33dCv2i/m3PDJVHK1utGxhHV2PofqLdjkjoR/TuS
mclS6P0TQLYX9dLFh/ZpvcUpXWc6OuqC/UIl1Q2Zr3iTzCrAx80PZVOE82eussxEq52xE5wKNMfa
iXukBsPW0hSwlu3cBwYgmLxhu83rKMzm71WGtmJ838p3WYA4aGe01SY80e9YTquqrqZ5K1p7qReS
NWnX95DIPoGPE19qRuW8CDV4IzA4clEi6718x5OequK9vGBblPaEsBE5AwaPc23c0zEqpO8UQXnl
KXLdRhy7WeBrcZM1rDqknJtcrJNyMg2/gHJH6b5E0J64iCcZGjfkFdNUUhG2t4qA1c9mMiy8nsgE
0laOsEhmx5WDDcrgIAq59XTmf7W4nkZUE6lp2PAq0icr2jSduFgjDCkWQsm9ipsF3q9bWex3YyWA
4/8gFnzE47sk3UaulqmgZhraM2rhTWKoi+t8R24iJAI7thDvTR2H8eRD8y9TQcJL4Hfvv2F1W8yV
ZZ6cZrlBO54HrEceQTEJL/ogDKNNtU9kQTEukHZ2KTjRu6Cu8o5juTfPoYzGnsMrlYPyGWKhu38a
WS9id/z5URXUqX6bMG5+68BMGfvFA51G4AMi4aQNmZTO46LvwWFSkm7Zl/fIRN4bElKF22QeQSAn
+z2u+Hl+SWbqdDH/8tBbJcit+iTDnnop+5CRtLJVctNrAtGw/0Lg3a1bhs9zCINB2xjcmcxcnVYj
0g3oqp0xPrspK30WyxnUMi+hSZZcidi95DHiAI4cbdmUR+GaFmBSkHXqXzNJ/Q3f28hXhyVzs4Lv
4C7jTO0dt/Bm3ib800OAP921+EJBekjx0xQr2jGWkbB/VqV5yr1OfsdSxIrZK2j7kSjF1JaJy67I
AX9k5i9S27nVwO/g1Lq0W+7xD1Rnsrtdl5bWw7RUcgx+eei5nYaTQMni/r4gns1jsUhgPO9TwYLu
+KWeet0B1ejYR4ieliJS9C7oeCwhxgml4DnR73B8cXi5F6yFmT1NQ46+5fOBdKaT/o6iNy1WDHzv
kkReM21B4ieeALx7pjxaBeTvkcrZ4pYC99ZVHJHkbw/B4s0ELpy/RBAjzgeKBzPJI53Ikq8T+6ZV
2CqZWrU0Z9mrC2eiV/YeuJFn1rt3mFogolHWH6aaixoQbGcTPSUAsCzvDq3ZM1EWohpqgFM9jzkZ
qtHrBWTIO/ZN2OYbFGdJy69C49aGldpJ8LvJxm0OzzjYSwPRzI+ugHtuKEYxaY/TcvXR7716kiHJ
oQxmYSK3T0q1wFpbLPRtHL3Z5N5L3kW9B0k/JvF1t1fJpmfUzmxuJNGUZFv5VR4tLjbRG5jK96nF
TniWs1N8AAlg4SEGHkB8L9DtcbkVnyttCZQd2qBqoHN5pWYX7Yta+VWqeztxrWUgSohYn3Wo2T36
rojewnvqcTHaTRljoxxV2BJU19bS/CxlBTzCYqGuHdoufPZW4U1NoAJJkWXmM3iFUp0o8NxPD2TX
YRnWGp1pbCHY76B7UPRHf8ChtQjTRasTi2n0ocNGVpgZMaRcTRNsUXFAWQlGJ8jsAcPvyoMLx89g
6Z54V2MDomAKqGuxu+2/cFIjBSUolopIsMRDDZPllMaz4wLd5NfmCXEupaE0bfpEHpDHsa14EC3H
CkNxXBdqYX4wkrc3z8SCZbScuauVB9Unl+2HuknnYu43RXxrtTLLymy20z8mFoiJ4Dkqy7R62zxl
dkppXuVDTdUUrBqELiAWnCmtCj4g+59i1jVS5T/VfvZh/TWYjT50bM9sQaFcIlN2nyM7d7lyC5hL
ex3U9krrLoMCbdAp2IcEbYjGnpfRX8noh5DcU2wzV35oH7gL5d71HLlYupBaj/nJ1v9h5jWrjLpL
VQrmUDAsPwEVomnncdSOjMOzgai9Svnx/pC3xFlY0bTF6opo6ELsuFYsszi+jiWDHV9pQhgRiuMF
fVLNUo05CgcZ1Wc1nynvxkDpKDB94hezmLysOE7VJKYWv5qeryD4piB4zJrN2EWFnMi178dGfR5N
cIg1CJkyFTfZW3JEx4TzoAPJoy3uCqLMVHi1C2+vLVeu6KF4j0Um8DqXndfPcFzsksfnSgLLQL0b
uzjEeJhxHudu7Hq1dmHuWz6ZxZ5hKTd1zNytSklQD+Dx46W75TbMywbOn/li7VHijL5i/fq30/AW
6Vcfie43L7AF2bqpTqADeL9v/t5dAjxBnU2nLQYzcF8snoTsD6saYSVBAOgjd2wFqYF8M04W/wmJ
m71U+WXW8sYjwwZ3G0mTJroN+PJMjR8SjQaLXE4QVCb0Xa+STCElCFwSndz0nbur2ok2lum4Ud9Q
1lPU30BzVLhtuc+Z8KmrE7Vpwf/LFAOJ/4p5nYYdHTIwjTPkgWl2yP57gSMVijKD9Qy+YMtPz0MG
Gd/j/fmFlaL0EL8R5MfJL/+ZLYDue3ESrj9Kr/xaGU2yXcxkw9VzfKpGr4Xz2pbEWCjnCNrQQo4t
TH2qkenGtwrXR0v39Xj2qwn6IhKGgKodxrxzrcJMjc6/TzyYZ9k+yKvshEqtk8h1nJ2BRu7lrmo0
/JdH5nUy9cDvObqfWNdVSi1oboEsKFTKg7wjA0PMMYB8LUopTp3w0RvyQE5lFkS0ZfE/TuFT3Abw
7QVS4dqrqlxJGEVHbh69tGOH/EcB8ny5aHasANWYLU5Hc0scjq8MbHC/mT7WoNMLpSMGAffo/N5d
ozlRH3cANnlNJm66T+DXoxdQ9k547+M5s+zjs2NqgQwENyCCw4laX5JMQrnlN0xJNnGs03u5M17E
DknqA3A4GnBKPOZDTdSHUn0bMk5wb//m2xMV77kNO2DR4ZYids2zckj6LdKwIpYKIMnunKh4kwqW
dLIKWcNKMC2D/7HAWST4TIRI7H6eKYWxpQd8ulmoj8xa7Vyg59/pB5IPFjW5RKg4VE6ruKLlohiS
IDtus8zap6mr3+oYG0N6WOrfmWRExDvPgZ1nECNbEM+yvqAiKL7qk9VIj7dXMK85U7odLGuSUt8x
cbOy0POP29erj55iAjm/MT+ct2PMUQqNMXZs3RXYMi7/C/wm30qmgIuFwMKKP+IXI6q6FmiSg24k
dGQc5JPrZAF2lFft73tZEk9EAo2aBcM3nJ38XFj+RXDbh0l0ViY7l8ultmDljw59Iv25GjR8Dqyz
Jp1QoRpGV+/0wx/4sZ6geqQA3kWEsieh086yudaddBVHdUdRpn/kp/zHImyISPy0cyZ9zmFN9H6C
4wtjOYVeQ/ea0HFFB529RVjzrhEnMjm0VOhHe/J9zYuFzeuiriiB8REt5DJ9DFKI3e94+Qv9LuYA
OUj9VGA5cjzOLTndFJ0Aq3/2DerifRrp147MhVHzF7V+0+cKEj2+CwExabausdHfpz8r9Ulaw389
7aDd1zQUTksVORLahmDSkzFnSO0GpjTgljJds63WiRgdOUobEv75hRxNn3kb1SJm+ZBpsTBt4zBu
r9diXjDvLk2xy2DITtbTPDFOLd/navd0d79oF/bOJsnOEKsJm8+Fqx4+HhyDIz2cyCT7pnP12oZd
wJ2LcK5CVZ9O7CJsJB8G34EnPNvXYVrigNhm1diW1h6MGQ2XW3u6vo4y6R3r98xZ3k+6S4dXsv3x
PC8IcYcmANtpxT7m68K5GJOCAtUlethSekMq83UORQZcNnBH1IfsjJmU7L6RIIC0Tj/Nwtqx3qFO
lyporHWs2WVy+afyi9O4QLX3dGeSkXiPxrUVMLmCTF8wavsUsJt66PblCSTJ+VuPE9CF+GBTlir7
ZCqBRaxJ3D9q/U9YKNroz5BWdar+qmGFZH9xQ7899AUL9x4IFBsj2l4xc0FwQJ+dX52kKEbkIReb
Tv2jjkcI6vTMWrC7/CwQaimkUpXdn1FyXx0PAIBpN57EkmVcVuMJY2DlDcgfUIEDykmJ17EB/0fU
u0StK/XYPplKA9lGQTRVhyXaR11WRomYMAIgUkHt2Z0WG7qytzm6gDA2KC+PnN0K48XnuJzMb+jE
qUAi021Q1q4YozzJfQD+iOiEad4P/xZpsJ2jeiJzwaf5DjlWTV+4LpgQQFqkID616SckYPTgH25O
0xxrFcgC95rhsUciURaxVm15k4yssFuZqA7Fm8LpsSWKMekZOr9X4K6nNnek57oHN3TcytZM+uSF
VUct2mfuDZw2e3OrO5I7ubAPC+wMAOq4AndsVnlCh+VoQZ2PxKLzBfJ9qkwirA41j19PlH1WrV6U
coDGPmVPmpwcxsOYwjZCuVj3WizwD7LxB96JesEykRdWZ4rZKWm796B/zdnpzmPHEBs/+lDzVlP8
wM9/MclNIvs+1N0eoCahAgmzuUee8vuL32X1Y41LQgyx7KLcAFGFardckhAx69DrQXZN7fXhS55v
f+yNKDj2ESUgWeJJOOexf3BJu7tFBhElfRpMGuelvHQHVSFKPlRVFkI2QbZw5pEBxovF5Ynatppi
ipy/8kWEtIiHUvCtQKKH96OMMgmK51e1VC1r8CmNP6l+J4gcxL6MzUpsP+pPTUkJvJ3L/MfgVXWr
Bob4bo+g/eUbqUYBnQKoVviDcYKomu/7ysSYqoV6ODsBtw5qq8HTG1DcrqP8t9sJkf2a2k9hWfhd
4nKhkkS5QRW7ZCt/8Z3Qz5kZQQ52Vj7Bk5oObxrYySJrOuUZ/u0NVSWmZAt8bQYNzeJvBkn+qKhE
tNpy+yHtReJzOIVa3h1vuHUzcKAkmKwDEs8dC6GyaD50DSlN2Rkblg89WFKkEvcDOGYoU9/B5MmU
owf/jAA5WQFKhqWASzQ9M/CfpL+Pmd2/qU7wMMDUNnEaZM7tT4Xj4fmO4XaReU5SF00C7X+MOUQz
9QxMvDOTBODvWKEMkD+G6aSzRIHNc5vXswQT1dntNDVKBJqb6yAvqym0h2HU3PudSholq0h6PDTt
XU91omJ/Rw6JWh73KBGOKsYGSWDUrEqGjVrfhsl6VrJWkA2mb/m/Et4KfsFBUCfTNIas17MY23rU
/h/lWWAQuWoDagsDp8+nTZBxbnesJFXRF1nOcdpclBm//dNMvu1EhFb56J9BbRTNxUmmx6SQ5Dmm
C7Qx3RByNo7W8gMey39qJ36vSYa+x8BxDTEWruBsEk8jhBxtSqBDmReVWTFMdRvtAh1YS+zm6DbH
dtLf3m3ViVNyJihDWs77xT7yn+jsV14kWz3yCvWaZlD6Nz3yFCtzqsXlKu8tqSGPRtDNJHOy+0Tk
fWCHj9p6etjVbASOy3RT12w2wqIkkEXTCUaSLamg5kxTTfnK8FIQDbUPQD26Og6r+/B8n0NHww3H
tQFq4LaJgpI79QK7U4JVx638U8bZNAhDlh7+kRKTaevjV+3CHAaDkx8nPys4VEg1RUPekk+PdxNU
6vQnEOItNRZK8bTj2aGqDtwJgpVFC88PYoRB+XnN8RT7KDdm2lcrBnC1fmMcoCdm6GXKBJjqV9xL
8ZbtplBZadKPDU03UXpeTonw6T8j7sUxBR5Zb/HTDBxUUJo2F35EVLcYxpT7aIJUq33aiww1dY8z
UlOq5ZYgg6zj49H3uE5z6Bcwn4ANdLJGK4Ey6bmkZiIr21TPKhRQCs/449rgvi2F49gxKwJzQ7xY
mNLwVR/EqFsR+/zPL4YYHk/emc2BUS5BmGoeDmSBGwAQxizghS/LeYpr4ga/q7NvptRmxmwb9vEp
qmKlcmwNUSKtTlf1WmYeB1PYdCyB4roLcfu5ouXJkllc6X/ZBQpUPUZg56G1uL0YLWhps42RZEun
3s5fAInnVzNUrj51dJ/DFM55W7Y3u9uPNrNqNxgjg1P9aygjMD6yP33zU933VrLXWUzdjLINAJGG
5IMf0VDeBI0WOgHZKGHKu4qy4dKJM/4FybBTCgveBrW1piGFHfQWuJMqaphGIoR2fCGehrOqvA8v
K8fnlj4M8v/V8KFBlqUE8CoXSOOy+xLGnkUG2kASN4btj44HNoNLqw3XhnAJ33OOgJ1Mc9cxRms1
7k5rUPQRLbyDG5F73TNqoFIdJsorbXAO0sh+dr1RGTjj7oNFPss/pXY808oNgL9LJTtB0TMDJ8e5
GfY1FfFXPw6e/AUo+QjxKUG2CLEbk5LJT2LTkSiqke3ZZpUHDT3fnKY6x+wT3i7R9cb5dKCaMkTt
Ty7rUHaHDQGG4sKgZTe0AGid1+6uGfuPMFdnlwjYW12ajeHXkQcWH63rQ9ruUdBLA0W2kTnRLuT/
f9ho+bm/MpOg2v5skNfxQ1maqJMvPnaurVxFAEYZN82cPJbFvlGHtbQp7c3kTS4gr58wr7hDeAfP
ZOsxWevBnFdnpCipq55hr1VrE5bzwtXkZ2akKPBIylcbOtLuztZdFZc8tmROKjiDCso5642uQ0C6
MQDDHPdO1k8/jvqfhTNUOL8sDwICd1QwhVxvyOYZuqzeyrpulGJ+/1xTEqa41lEifKWW54QNaR6t
lz17qneWhxsNITcRszJ9Knkx5Yvbr+eI+SumGpEiEpOrM+uS18TrCUl+LGK8egpRvGE4c/UfxohM
rhhxqou1Lf7NdHX1f5pFBWe8sHCm+aduZb9QfE8rxJWYbDopRmReSqfsUZY2JscbjJuUxef5D6ye
+HLKSPwQswkT/FErOBmZj+eoWRfFIO22lpHOMy2z02U6cN1YPSJJ4pO+g4lxkmjwV9HesJe5qYWY
GjwYU8Qpj1ORgl3nLjTWpc120ksNlFNnfqTsa5DboOLGxg2TC3g08nB2DNnCWLHQwkge9CSruLfT
42sDMPyxVhtm9tsXuZcrEEVPtPoF+8s8InHQnQhXNzUfJi/QlFPSKLc1wMHTJYoStjrPi8oquJGk
UqxR1+s0P+dHjyN97tDNMSEfzSlm1mfqHj+HENg1CIs+zJZz4QSQSjvukP7ZXXXyyAtHlexWXeRG
4q9WoSrTkr3mOJ9hZkolTS8ywID6jLJnQV6eMXAesVQyyyqxCXmpx9RT5zmzk0r6QMQoNiFgcQ4Z
HwhV5vwEaa625WLEKRAccSowiacvXA1NyEhwsLCtCcIzb08sn4a8FRrnfVxKuOj7BV9oKHD6fidb
PCTVUgJDuP9U47kYLj5+O+mahkX0dUZ3n8MJcGKUMF0oyJeS2Sj/Fl216lyrIAWtY7tLD9oxceRj
gilCj0bU+aFpZoa2D+L1xTzarFtYioWyMNykeadtC79e0q8hGIOasYaQ2X92nHX+a3iPgLta/sUh
ySLoJo0fWmxIi/OEQjr8J0lhxdr41dkK0dBdddpGQ3z8eh+omOmel23CsgLyRg/+qxLT6nVqJjE0
cUqAOdgV7w0l0ITAac9TvOFjnsKtkEdDsHzmXWU+uV3VmxCyHiBdOe3EVgRhW2rCnLHmrOgHGqia
W1ErS2VWiybeUfPrenzK9Goq53BkOtlMDAA2bsf3GSK8YOrd5Ep7wSsABXuWFiUTRGWA4fMqNoM1
J4eIzhAMLeXNEe57uBFUEAKdA+VdYTJHDPQJLOQsEzYTgulPTM2FrAuOlTuKerQ5D+xKIfS/gAQE
w5BUnyBvjCHECYkLmJLu6ipRkF+NN5otBcA+jDOnjVa03MG/Kvcdn9nfT0FRTClgba4YCgxz8+gd
Gzhkk2Fw8ILPFTjyOfo1/8Rvwx//5hHZFmTqZ4bJc2wKiwTJVi+aaaOakxTWclknwtqhVtMcnA3a
uvGAWzGaySgcCNlGayzWpJLJpqEMiCf/hULRjTgHc1dqWQqZtb9afLu4niCtQ92kAu6TR4SxJSZS
f3KEV9Wf3JOn3l/b+VLH3H+nzY5kYDz0lIluwQyW/6J6CxR9i7gT1E7mrso6P0o7yaaJ261jweur
wzO+q19nInbcMFXbWO5hq0QmO839sPwNc6p/CwUSbMp6nmz/r27+RWneK8eyEdesX9OLnLJAyRFV
pkRZwEq7eOYz48LIZ7IC5bxiYyUKjJlUGXqJxjC3w6ZyrPmz/7Nz57TI1U7I+OLARvVQUyAVT+GF
RTAmHvffcHUKiRY8Y502WjnK/4yzEpqF/Vs9xJB9RYQJdgDQxlMmD5QZqt17DdeF5k7QtbPHSS6P
ZRYV9dmu+RYIf3fJcLh+hxRclut9dW/AKcCnwVhcnfceM9aqMZM2fSDo8a0HeBG2icUGrViulMkq
HSrE7CzWRxXkZWx/dbwr6XJlwdELJIHiZAdMNNec0msXvuvAFcgoPb5OBMae0BwPV0QpHtsuvZsv
wXvppQ33LdqDNd7f/3/R3D7f2CAYPiG0ycTh6f/+v4fLQXN+A/wQ/YKIOAPCCkqxRsnpu3SprbLZ
yh3OppQgtwNJkh4N8DgW3GoiY3KzGD2eWcGgX3Dtq84waMMyVcRLvYZoWm3C5e4kWV36xf2Y9v7+
/FnXAtY2zgI0957yR2riGyrgtb25z4SvFUhUYioP74//yPzSpIP897K+RbRuwMlI/cZvE3N2N51D
MLimjVibPY/tFmC78/dHwzK6BBo7kC81nA86E1NWvXiqYC2Hl/MtcJ8afoG5TfnCIb9DtdmlYkNG
3Zh9dtfGz+QehEqz5jj93z8O/1ppUoUxDvp+GUNoqgiddkP2zr5o2GDF2/edm4idxtYIQDDi2//4
CzPINS/reYbu2d2sUN+Uv7cO7f2YmaVd3uMqDmLHV9Q35mTrHjp39lYJ9d1Yjkfgz2qhrhlBmWIX
YfvC+2dfCYi3rdQz6lBgO0KbwWpcA+jrTvLDeen6NFLlGeDW9bC3IKeH6Y+Uz3/J+LMEa0RPlTSy
4O3Yr7VdrClOw3MlfXdYsh5m4UO6FiEkn9nodV4xcsG93TKvK7nR/cbCE8+vFJipCTRfRzF8dpFt
KH8RN4UIiOpUueXjvnuhqm9BlGsaVgjCOmR+H9dDbYrrbirVcxlP2LFhNkNd/nBVvkmy0ZPDFl46
ZkyLG0Sah5FSOV3/ztJyVokQmeiKabSD6eUHnB35SuFBZTx9pXcAh/wiavEys26Pppep3t2hGMUY
2XYKq8Na9j14yASe3EE6SzMpzSsKp5bAiIsiJYjCOMMmmQjzsTnmhTnJ271titkdbhG5YqXXTYNc
I0xQH8zHq+hVg+IsbHEwWU2oq4gnKD0XtjGbUaOQePBfs6v9SthXTjt76U2d97nMV6HBTjelhb5J
+OK9aEXpKCWerHCTRSdsui4OISZNAMlxZ1DbV6XM7B3LPY83MNAvC0TyFMtLzbvZv0nu3WRbTrI/
q7rHtO785lbjH8ScubzrqnD3cOkJ8LUjKNAyxjjkYwNEYbkP+Fnt+8FkxK9hgaI9O6Wk6RVNXzfv
K44PQU4oyZ5uWdmZuPlAsnB5j9dNGW9EsWp5tIYNfb0kuFgqWxExzxndjjAU7JvrrhJ+Uh8rPM1a
6xRm5R14oP5J/utAVtmjYoqMHMg0aNdYmq+L6/AjmaFxSle9qDlIy4DIjp5a6cY4IvefkpSmpMna
pkFsOa8Xx2FZmAv076wOp4kdHeAWST7YtIq554Xqite/vMOxmxLKXA618tS8WuHFGrpooM55LDtq
mN9cnWLl2sHn4kLdo+rvp0pE20yn8qYXZMQ9xHJtgvtg4vz0g586g+ZUyJJpm1k4Y5a1v0nG7eWb
cDrMoonAbw2hNPgcJNiRXiKXRXHsdeuD4vOHddn85KM8o6O6Z50qLdPnuQAT84c/NGR3H0Je2cZ8
h+SiUD2sxmmWzEp43B7rwOBSyYkVqwBbtqTPve0470DH96kIA8P6//C0oZut2FpofrlJOra9fksY
MpkzHkOwK2zCX0IOBHMcKDBpq/QnALqkRHjRHCwRVUQgGaiqf3p2fPJjUdfrPxFeW8J7vC6q3ktd
UDF5h7AAkH4Vd+IlkJv7AtR36CRvJ+m5QCXWj/FtstAsQUXvHyOXslOivh8tmP+lJDiS75tEJJDa
+ZtFrUiAmntb/8EU1WVbRIi953D0nD7TLUdUP4gFtQLqcy2v+pqcWNR5oGpoDlFJPnEF5KjWgEZf
jIQrX87HWG3D412g6VUfiV/3msa2jGwc00+2t3iRfDc7WOOK2Df96vxPknbJM85bMsxXTGg62Evc
fzm6qMCPc/kNjjqG/htbGw6tlFwYVMefGQzZbtx/gF5MKs5jyCBVEMXncGfQKd4dAT+juCUm46cC
nqubsM3Mecc/tmM5bOrqWxs6TB9VlZo90VpNW2pgTdnqVekiZnaQ5cOSnOqQYyY3SxivgKHnPbxJ
SdM6of6DlOlFttrhO0amHeUU+D/LDzvcXnuVAYkrSW3Dk+91eoCPPKIC0B1Y9ejX67zxujRLg/77
80TjQ6bQ0TrarJEkDhRne5k7eDov0je8387NfRNg6o6Uw5iZ1yKvNeuEB37SnMNSg/526Dv2IHSK
nBpbOvH4+2Vy2vTOk7y95qLZ0ZKTBnVwsfA9mmV7M3aZEZc9f4+YzewmLFlKl3XlS58/vEAkzUFT
aRkjUc7Ip55hWgUQz2JImwWZUTf1tWc5a6oblzDhuNfrxs0nQSUN0mEEMstPQV2/n7IcL0ws0nTW
dy8oIVe52ADKwWB8rMDT9OoJtkvWvyYPMdjEj9eP0mlmsoMSyEqFZhVGi6zSuyjvBqbvce1CU1H8
iHLPMHgFysaFIbTWQHRAx4e734fLJvD6HAcWB94yAvKtYMWpbHMXd8z2S50XGySjVT093a4rsvlU
yPHGleZ71G4ybhLYxC/umAcilVxTikjpAXiIPBymfJixyzGKc3uK8gKHYMV4DhWyGAtDHb5zQXFR
e6bEz027WUp33GtS4qBd5VxgcH4ovjn3gNC3hsS8cdwkNl1af4ZlolD96Ou7XMRY4jK4ekLPuopQ
U4rExCET3iQ6XRWxlY99LZ8pJBdktqGrOslym/IuUFGPeGP8IDO2guFSHfpyyTrUqmwA6ZE76RSp
BKsQCEu7gfSUCZJ1pNsZQAPZyLEQEszYw2Doe+DpPOq1Yz6bLbSTtPgcuQC4WiDcE3CHPV+qgmoO
elmZCS+OiTi+EQnbGbP3UCq+UyikdGzFcY6uThIoXWpjHDLKAabtjFqQ3G+v4yPLSVuKPA/eWJkp
llvJdjGIrJaUhWwQxcbAbloyIxutCMwFMmzuALSB9GMB/JCs5X95q50uCeCatl44bZ2TculDmlHy
EWH+QKg7xyZzRg/qbJkbm6KF3P8uJtm3h9MCwIiJbwIkul0LWKrVYYiGtf4H4bl/6mBqUxaeucPI
pqYHicylFjGg1YQdT8tJzdFZVhWr8jpFdGS0ouKNPhZI3a4WJmObKv8PYvg2oa9OWNq3Bu9MawWu
ZoHz+MP2khoJrp4gqLgXZ9s1Z6ACkdQYUKUQRhscuQqoAxJww5kN2sK3gO13ThRvxheiyGG4d23d
smBqnL1vg4b0+pgMFS3wmg9eyyEo4CjqFvm9CeAdegcwQjgoq7qgx5mnLz0l5CV+kKp47vRQyCHu
1CA/occU5l3tz+AHIWI3wNUyIXolNrePOJ5vO9A2PBbUniYfsrKOPfzRutTEBHQZuo5aN88ee0wP
vCpnKo3pDXQTzWLUrVclYNeMx6X8fqeCyBPiKEjt/Eq9LmakqFlTznwIfJfDFXjyEljH+euhHdSw
SrLUjuhCS+gN0Bq3y93pLcfRINoe6QbiW4CryivYRF4opdYGzPDZRaGITuWSNMxcnJtF1193P/Nf
h+v0aAP9QBp+n5YF9lCcZx+uEH77+4ISHmP/ITubjNtvmXcL0U7WsERAk6dODhqHWAF7m/hzC1Sp
b2NnZXkEZL764cqs139clt3ZkukEO8+zI68SLu171AhbYYs3cCGWjnY/rtsGh6OFaDrAcqDJo7Q4
ljB40PSRxJhmUMjirahIrqXloj+Hg+fOx/fjXPKUWazMO4zUap/euhJREiL0HkxsOgtmWdqcm3d4
e/+mYBRqpL8K3EcAdkHUvFv/l3OC+SK4kEnCO+XnaSgnNuTeJvQgX4UnJhbb1cFK00iAgn/3hZoD
KGqaII7kiQs4CIAmOaK3RpzdjDay8lElu6U6KVd61wbTb1h6f8F6tkfYlmDXNE6eXagRuR424K8D
bS7rtzIvph8L2mpIi+C3VzeY0xBX45intc3wteQkaSHWpsPtoQQ1U8joI8RtfuiFe7s7um8/3jL8
cbihawCeow8TksxFXgIlcUrsyq4LxYU5D5SiKbvTMhB/occTvKucdV5Ka3GUYXhcFtRQOZmViGrg
d8FDHRsmNWzDhsJoeupq+2yuhcTSUtQPvEXCR43r/ANz3YM8cyHaON3roOoK9dSnnRA3/bFb7LGW
thcfqSRoAbF/11GXPKErIeeuznw9oX80MSXJsGo7HZp+YYbNTeGwP+C8t7WgcsN5J/ELa/UdbIfw
cAbhNtNHOxmdAuAjaTtX/Jfco5CZSv8LG9JsX2nM/bHELGTFwtZg4mzjLelbFJ8v7nGuZPHWLxbb
ebtmERJ54YY7UQP/CJGzcJUqd+O3sZr09sefk+w8DImT3G2i/KEiCgVwT77Z/oZJC4zPvfrkgPnI
sTIMFukTgCAEgKef8Ff/HajWfBwDp3cUlb13Mb4H8yOdxApwGBQm4gm9DgTIgbjUhhUsS61PkQ1w
wjiNDTps9aLKFk3p7642sXQpG/5BHoe4FapdQ1c+taYQ3FcnaxHuhaU2kG3lMBfZghW5YEQ5AkZO
RCT39arrVpM2WKxRIkC1d0/TE13L5ircrbwiN+k5mvKQuwPpJqyFytwtfkdLMuhsct3+AOWT+VMC
ktr08DGcYURbVKFQk0RKIMxXOlu0h0U3KEpxB3mX4lWaepnYQiyXhtPQvo2Sp1V7QB/8hSPX52eY
pBun4EAfBLUChzcm7STHZN32ZUkH7V3Xy788398EBTR9IS+qhb0+b3fVERY3h/Z+iX1nuGxNJPCq
OrIyCMnEzezUnP8t8oAfl4Uuhb//oeuT3GwdNUQs0qt8+D9IALZe2bngSIIY9nSokZmx0n+2REe2
oH2mgV06JDG7rcR93bSB4Jrl5Kb8mNs8kXHXiUKMHfBb4rx0C7OirnGMUsy7PTRKiDqwfYb00lYR
WF+ULuOWIZiIEJUVpu8QZtgovrsy5xyhj9KcbIjwFMMAAm4sD6eQ7RJkvGs2YtBlunZ7bFxPZ//4
tzELHH8XGvVqHmoIzu6lZ2Xt6RFumpfBUzeGMVBhaHKU7hh3J74yH6Pdr/7xMwrjcnVscDOO2vhQ
hD4cv7mFSiIQ0yP0SRhYglAn6B5nhqrrtsJO4aaAn0PlaGKDgdhEiBVWJYe48otyAqKJ4zDGFAp8
jBqTv5ryBX68XBUuwyUDM12V/PDb7Ofpc1SPvWMCoCRDr9k/mG3UBzVfgQY8oE7914UKvFusVUfv
UCoM7nai6ldOATwD5AipWIXXc/1O7gDWeqj9Vfa+O8X7011QA69L4zxjLCPUx0a5u3UmfAJugf1z
k+0NGqF6aVk4vxlvJUSmB9bNkV+HCXJJTv/2ryPRBj38Axv4l4OvYC1OVT71+83s0omk+XvkPLK3
G6Y9Jj1jcTcM5C0x8QuK+vYbC+IgQCRosAymffD2cSDdv9WZArUjdLDyIjvewCehdbJLp8IdCKux
/TKsTBSoLfx9I9HAFKeJsDZhS5yJZcK1B78C0bPXTREq4SmIv/ZZelf9dlyzVDg7BK7r2bFmD/OQ
mERYp5mGCMdPquRBl8ykw8jNMOGChjqQBOvUSNBaAYUtN0n//IpYWzMefQjQrWpWOp+DrTL76D7z
NpxHwVdiaupL5Ml2TTW7OU/xubkL7Qa3Tzzchp2iZhRClzn/0IE1VKqwBpyd/AD1M9Jejb74dbBt
lfC7kN5hXs07QRHKmcOjPmhzgYXrh9AUiE1oQZaV4TRizIsMmRGGszn3BpG/79JjIKtwEOKhVilX
c750mndTOTKCrbjww0tdgtorGSVQCyT1egIUUVLApUPVIfJq/0hTzjHPLUgahWCCYIkyarDu9dVf
gYYrkqOu2bYqeyLiEowObC5afOZ8h6r90mCxngEAUL3ucyXc538G0z/YolPhmMQEJN2QNwNjSMp5
ojrMMlMdTY2ZqJbb/iNrECVwRsAHaO9GiRe0VWk9otNmUqxXzPCoXVJJTKbxB310nwjaGbnJQ5BD
fu7yVITLdl8mRU/os/GHylCpH8fDWN8ldKR3BuQ5oT1CneiI646NngrYPHd6+/w7L6KiizlaitYG
ptbR+I0OtRK0iTP2FtAIeAVcNo/jX4bmLRl8S3Hga+SdiTBGcReKm3ZxsHsAP2b3bCWPWIn7UWn2
pIAh3HSG2+ED0z4oTAFMkc7TZQZhbVyf9gSeKNQ2HAN5IjrhR6xSVvHxZ15CafvW+uuPRy9CVCjc
Jfa/GssECIWRLu+XwIJiewqHcORYb1YM/QZ4PgnzJEZtbAWdjwMBUAmxQ6hAImz8asttt4HmfE8h
eC64XAVBTHm2WS5TCQ8Yq7TLl6GcB8MY/DJ+Gvipz8bne69KAMg520dusxUmN/RRkmyLO5PORzL4
E6sbI5te5l4+NrzaFSvjk4QeGgPu6XhAqh/ODmzQLMC9jvb6GWv3F4D3jj/6BJPZTQDEePStROV1
JoEsNclhM7hP7YE8QMpvZEFO/ZkGK3wW4oAfgCNNhHmWXeNo5drrzJCiB4JVZpaGX+EhDF3y+vUh
/z3fL5xQRkmgJ4rpbXZK8KrChToe4fgf6c0wITqSW8q7PrmAuOU3htEa58GuoOmzc/8uEOGXPZDH
jWiE4uFLNMNh1kzW7u/62fg0YwNwicH5Icp/vOV3DKom48Z4p9lH5KIa3G5b9oTiMNaPBMk9s62f
er9U3xR8O80o/2t1SQAXBBp/27FHWwpF7BM/KFxaflSMG7GrmHi7JGk53qrRhteB7kuMg/t5/vjZ
wPDaRUf1kYPwRv7coiC1sgw4CL2v/GOzmiIQxFOif/F7VnpWmVFsBOlPsKTAtpQaEy7mYnso5YTI
/YboZ+J2GSsOjUX20iaVTatXvE2/1VmnZyFT7Q+BMhsp2OqgdQZCLQ4pMxEuUp1PKzfxPfTiCrTX
XBNhVuo4+KzsiH30q2D4PlpH+MfWVMlxGeKBfdufLWDRjVJQUArzKsp4HwR5N/T4OJlcxwScDsjL
TsVD7aDkydpjf8sU24OHYZJH4rQ+DfHYGFqy7YX62DsZAOpbWXPB7QBGFXByKsYf3nds8Nr2vxaw
INKnwVdapI8RGIN/ZIrI3K26Ur6MATUq3KxCNgFe4crvnjUGiI8iLFfyKKljMy7DYlIFfQ1oZDX9
JOKmzhpxboXx61P2ukxf5Kh9fOAVmCQjbSn7wvqRrvMy7W94uoXSn0ktF4Nvcgk9ERacJDpVnMtA
rCrkiB+QgqNapm1Glo3w/dJTqWADRPfwVlWPIuYr9G9Bh/9tike4ypYZuY4bAJ+5ksusV2Njpi6K
hBeFfl90wKOjQt/v9eVZHyYO4FMRVozyigHiz/1AmZTo0h6Z8sOnJl8UmkfqrRf60G8Jvn/bEUXP
zw7i4AQXwsAr+XcCSyTZzyfhPeZyndgNVMpPbHAHpaNzsTiv7MC1i8Jznshcnrh63n+MvsTg2CzD
Zo7AcGaJnqpEACZIyv1YR3XBKVdsghuVFekXml20akNsHBlx3BTrdWUpz44eUph/Oo28hD34AJV7
JviAwtGGH1ATctpRLcKYE7cNuI3FGtNvwEE3p1C9tINAFHUcN+04miadE7H5indNtB6ybcKPwTXc
KBgBl/lX40LfuxN+rl//TZgPSRH3P/qEIV7ha+ZRSH913E8ZwrCs8xHXHFVuE3NBKwZsvMOCi6En
8Ug9V+ZuLO0VHITo27g/6ShDux8mDufRko3aq3SWM8FHHqKG9bR5Gal3Pi4Tc15v5UfSFXQUtpy1
Zn/kv3JPsH5xBaI/Fcrl5y2GCSFBb8K7SsHH3ydzBR4YAXlcj8MN6ONvZtPQkTOrgMbUXXnh3L9Q
PMVftk6yfUOtx3oTMV4YXxJZVukDHQd7dONwpacRcLKcdaQWK6AYwqHBCG1UGcktJ20AqHkiOc1Z
4bPZBEkE+Kqcn5GQmwPZcb6rka5ZyCufswrdj7uSZ3YvxrrX7LJynRzZJCXBysk5Q9pQdP3VMPrW
ZlBQf8MNSHckyhtNhLqg7//56kffJnaeATpn9xhHLzTuxtwDOQHyDtBLbzteCVlSgn0n/q+qbd/i
vSug2sGaAdEboJk8ovl5jxBZtLkU6Ah3bQ9A2BLa0FJnyTtm0p9/sFT4FqwMWay4r6F74gcygLuo
K22j+nKi8XP1WF4wq53il+9Azj4c8gmGkQIyVY8giRGSwxEzSFdl2PWCUXKf3XvVYYRoRSCHkq46
hPaPTRTzEB6jx6MZ76Eo4XNhcbGEQJVXZgYBok+aZcIzOahRedoW62lrgKHzbx+V03+XGrjNjlwH
A99sHgVKXpbBg4qLGYthbjPPhVPm2Q6qhkTBYmpG9qU4OJUB7LyIHdS5k5rYKfTqdvptZZb3KcAO
EAom1CvKXXvoDebv3rwm9mS1ITi+5Wtfj4syKYf5w1WAXQpurfiFqu2nQLJ435Ag3SrMlLKAdj+b
oXp9coPu3lrnZYfIDqq/wm1Qu4F75EXXOJvkDnfDyBGA30sRuprN1Kjh4HL5AEGndjm1Ys6D6LGN
t7bE1xlNKfu8E0tNVIk5Qlt+KkYBx42IDd3bGcp8HtcP3s18N5G2RrVqOjoJ8A6o0jt+KarQ8vAZ
0wxtFjJPFhBVJmnPjvVZWXKAu3ulp4N2z9ktqL2GyrIUyx82CPQ0TtNolB1asp9SKBsnfUkwnJ4c
mRYFOPjYcqsWzREAkRrTjNwNa/vQ0Oo6Al52WGkEGr2uSUyOvxXoOVRXEg8t8FJP3XbVQXP7HaVp
89Tcp9t5mHugWs3WZ4YkP16lV6UFzhf7Yb7h7knqziGVRL3dzQU7LSSZ6658k8Cy/LnywwtXsEv2
l4qe6IK29kfHWY6VpgSLKoRjW/BDU68K9LnQmODYNU7ZHzqnS211rXeitaEUulXZdXm2f0oDCl8T
FMCsG/R2hB4U0gXgSTSIOcywRC+AdXD1B9Z81Y++aKL4OB6eXE7H6q+7W8Yxhkjhgd6af/ASrKPn
dRUX05hx7dhK1JxNiQklE9OW9jT/joSiB2C3NkzYqVUDy9Ar9+6eDu6XdzB1O5KiESamz6pSq9HI
2/ye2lFaFjhKAJ4Mg2+ZvEcAO1M7PBv0x2F86OKLX89RqRXhRMfTFtKdai3zE4GzUj5dafS1zMl+
YWHNW+nAhQ+7H2f/trBCPn48DcwAh6qv6o7Hgu56QevLOjyqrn33UJ5ffIZL81JRyqEL8j70ANdo
k8hek76qaVmuE91x+1GrlklSVYndE4l08fwQLMOvSYc1Tg6apTq/KGpm1GoPu7EjUOEBjH39yGDV
/+ggx5DF+D0QWXYVYw0eaGw39lIcfO6SsLHO9UORZfADjPQre/9EvIMqeFaicY1f+35sAfB0Nu+Z
Kkuw+S4SM64y2oFthxU77/ybQzKmJgkmnHZU7iu9rX6n0r3GV9MpxwZDI2+zID0a+t+1V/CU6L4E
gBeih6DdOfOVrkbCpWemIFjTrDbvKbXzYNe2t1gl5Uzdkwx5vScIrPqdOX1IG8YJ2Xm0rz0ZH9GA
vlOoZvEWzGwhkgTpCJp4ca5mHE+LOgN+JwYvx+TSoMTuUsggFb+WhVA/fvNyNXOScoF0k635vjEh
RvDzMFn7sVcsDVqAUZmqzm2DjQplu3MldrJT1yvpOnKCp7wMw8nARZrye6CApMV4ZShhjrk8VcMb
/mKIppmNnY00aQMR7OIJsf2VFtr5i6JpKdJTRXI2+BewyUYVY5DR3CXr5IAHcJ7rNnkQ2UUGTIJe
kcj/Hom9uOpcemvist0/h0Efr3we5bAruoOnW7QHNsKc+0FgDEnWx+Gy/I9Ufeo3WkEx1CIsTmso
TRQ5MMKwosKYqCWur9oKIn751Pu8ikbuGpctoAY1jfvMAV9kL4+ZAy1duTteN0qoAD2NL9dwDKZA
CExdkNKT4LCj/Tcy2nd7mPLsJPeN7lxOkXCKc1WfuQYYuTNCf22NfbFSvDPU5g6YlfL8UHaApCHI
AYHzhMHN6g6bpxJYMqNqiZIseQHsBE+MAcIsFNVTJpt4WKLpi0jfuFI1bso0f+iXU5Yuk93mTnEG
B3LZEGEzjJXj4VBMbnsJUGrGufoKR027zKLDzYFPc4T7Pv4yzVIRMo24EtO7E3Bw4nydA62BJjTb
osu5mOWVJWNilPq2GYBSkjtESA9trqeNlTs0i9kQY6eM7iOk3tnz9LFVHUXwJ3ezzfoTERtWXfGg
hndUy9g0uhbydz0s/FYMai+A9hzIo1tOhXVG7I8jntiprIs5QvINbtEz4XsKFNLT0EZqswhD3ix+
DWw2xrd8vOaKqFQ/OyTZ+LAYe+jW5+7hD9/30wNdXVlBY2BwGrl1MbI5uF5CsufTgH7Xzh5g8Rvy
44OrQNA8HbfbNDL1YNYtMNqxqnTNOiYCMz0raD0AchAqX+f4bznWkNdmWS9ypM9tgkGZUmii7wxe
LXw7UVI/Zf6hZ6qDFwPRPltU8m8YuaHrSXjP9EUUilGdskhdsyJuNaXQsJoF+ksaHWTUm+Y0cR6t
7X9/JffbTO40InrGZHpVrbkwER6PtFwP1cWo8lFql5bgNBRx0oeBzzElehE0rFMIciHdpDNyb5dt
kfGmyIXXc7MqcywcxPjtRenIMASrUAd4bMjdbw+qaTDbbDV9rQoVrYD6tggzuB6VEWAWQvfFnJpM
t8Js9ypDwZV10cJAQ2UxWUJeaTmGchFgDV8c6U2NT0hzkNFIs6qaEtKpYUGflgmFpEA6byMGgggt
1IH6hVFtRLMsdIUqpemnm4SVl6QApu8akmiX3DsInyGnpKhW00bklZEEvNcofgjNWJ41shyb+tT6
wdT0zK+t34RyhRcoxOTs+J2hU7x07K4ZLTOeJYuusf3AHXsQwKwYRks22Orlq9IlShnfBhn80UDl
PitAMJZHVN0GWrwNzwIFANDneL28lzthpBJHbmVqq0Kpkx9KnWBRFgTYTS0dpUOwoyn+LatM5Qzj
wP7xAE9ovCkpuo7PjhQFg6oUmUxn9LJqAsR3t4RxkcjaVsp4SQpyp/mChUWwYBiZMUy05/55HTNK
Qt9j8Dia+vUk/X5E0yO1sSLGGRUqwtunijDgWGbX9rgm2+Pcmc2i6xdYf9JJqLTj1wZdjZc65UaH
8LPiRPIfyRuPKWHlVylb3IbB9TQNT/VcvaUEgF+5YzLjmfjRAV1EK2VxHH1HJhyv+gWlaovU6+cl
YOIUcSN8mLKa6/oAldjddEcigZ42BZiWoZMTZg5vc+LgSbRwa6Va3pTB5oPqorqBVGxxFN0rZ8R/
NUdqt2ckIZb9aqQb09hZHKYoXvW8zxTv79e7OH/oCpLWg1SFK3suo2Sp9dcrMGdc2woa8xy+QbED
o2q7K7Ze0E+zJpnL0/N8njd+u1yB86Rf053j8Y3blrPSOev+KmvRKvsqu0UYRp3v0enVEJsGIU0m
zwS48+eacNRaGkyqraw6iHupDfeEKnA0iavkQwkD9f7r0c4wdwBikdY8MPUVy70/MIjjbnq4gk2I
XgHugrRo/3rGrtj0gXmnrJyXDHO+EtGAvTI/3h8/Kj/HSJ7NMCJyWEkJZz6ASNd4d9lkGe0b0hoc
uMVFnPb9UgWI/mBIkAIvRpjjLKwg57ZFAqpVY5hQoYkeBZFyK4VYVaTeAEmvUX1WT5SRy7mooY9T
vlf5H/hqo34YolbKpTLzYjGAYJkMp81Cz5csKNj1kvo6tSG6KGJkLwR3h48Ky3CA7n/OdHRXHFmg
nrw5evvhaqe050YqDiV7Zt4ERxb1Ka0aJABiz8/D3OLJW2eE0n7+yFcVzsUm45+lwOMgeWV4DvG4
leDKPrSIgORzNCeGy0BRTmL45zeVFcNI/wZ0JIlGTYMZ+MQaLwpqAcBnw0qZDOh/WNv85isACh50
YDnYWnKBX6cSTCIg76Ob9t/UPr3X36ZUezdIcFILb5DfiI7zMFR5d5pqm5Xh1gDEsM0jzbqCNnkx
rdiXaGNsuglJhNgY7LE8iaHPIo7/C3kp1UiCSxdz9i14b1erOOhnoIobhRQNVLq0vmDu4Wgi6z2Y
iH/ay6co6BVxiY7DsEPII4giIgGMFmnamUba4mVlbEDBQ4dE5sbQ4F3FDf14on67SKibATIf1TNO
R80mxyYMI887lKte1q0woeM3Ykpb/FBqpunhglDaleAFI7EjcRGZhG1mDUFn/sXvBRvqh62t/DgO
3lk1nZRea7d1/2VyM+cbsKEttYA0HvP0o6bIEegwhcdefblar8tYDVFU3WsMEaXS2Hfoto2rk+ms
IYIyTHQwyUdUNA6mtf5e38oB25qqSSwXKWXQS611EtVe/7Ll3+8mpJN/gdvkfWsQx0/HcXrQ7U+t
vIdlrVKCfXRkTUM2URc6m47m+zSC9d8doTb9lCBuT7HdXnGA0idefqtf7voYPX/pw8jUQ8N/DuXM
xv1de/sLpAyqSyEhUdb9eacPs74+xoIB3izCHSiGaGvB66CWs8bjEnCpcBdw2+SajR4SlJNFEul7
jPMf6F4A0ibkqFM1IF5m93BAK+889mo85EA1xq4sGM7vzfQ7c6P5+7+fzNZCGj/BgT8gOhkxBe4v
LelSkYts7eYEMH5+C+r/Z5TS9ZNcTTGWCC5slu/BUC/ufjal6np6IokpJNE/pO/rHP48Je5D1Ocj
expdWc98nIkY3BSMUBNNmR+gtaDVg9er2/nysWDQGxOImZnmo4DitIIqmxTaVSNtvFUlU82nrMWS
qfQ1lM+pXDxlJwEhPOJ+v7X3IflpHDrdYiaDcnkUk/Jaa42z1GByTyz0Bke0I5WdcTa2LNATje8c
btvVZAQp9HrsnT9qC8XRXG+E1ar902wRye1KvDA7Ek9BZaSQQ+b+7+wdwvsrikvquHQUkeh401ZS
hmJTGUI6szJHC3O1lqg4Fyr9ROSziu3aNTQkY9JSOhdgRlgA1TyYDNKACj7tySIkmWImYupKHeS2
vjREkMtHDk3Nyhm2lkshHtYQmBO0XU5LZx+Ss/MNPG3XTj9FM0E4A89lMriSaCkmcABVHw++ST5g
wByW0fDb46hKsOpdQDSR7FWXjeqSLlHKvl0bwTTI5RkMoPg2b3H3PlHnnh6pfsPS1B7zlqOX+7xk
VYjG9Mhp4xOEVK2JFgbVidXQ02ZKGcWs1R/ajxe12//1g7bzPdw5LhdePW9VGsT8TRJW49BFSWSB
OKInUy9Gqbw2epaIlIo0tKDBzGNyhbJGL/tRoE8myRM3SnlHVz2K8KRGpS6XmX3U8XtNQQUrOwWF
k0HiDiuJbUJtPde2QE4YNQP+dtyFqYg6ylEmLNps6s65ipRqYIr6QfZ+S4cwfR0JxeBYntT81Kci
3+IUf6I7C08fvX0d83Iym049jPCZaT+awfU9bvNXbPdkCdwkNTLqCuKiiXrg5+y2bBfPa7nLezeA
9MXY2nBqO35MnKdNyVzsVKre6pHv/5wTEhDm956X3m6NTlbJe39mj+aB3ltac1fjTbelA175HGnv
1xFe+PBu7a0Hy7cVSXlQUnbkkaL/4JzZio0mFWyXgQQlh5fBHYrvERLGm+iClTQ62gpIlZF4s6jo
t8JrvyhsmInI0I8wqfr8tzyl+OKotj1W9H4BHinu4sZyFh0+DrUChv0e13Pb0wV2mm+g91ytcG5Y
E2WH9aFyFh19OtCnkdeoy6IMTSI/kloYvwn0QxmhH7mwogiMDHcTREhepb5xK3pB1Mlh8vCk8p8f
+e/7+S/1ELTqdL9ukAYmA969TwlSVmnjljavQk9mScIJUW4QwdKp7DMtCMqYhdZSCFQ1qdL0NFWy
2L0ET5JUBYYKcxVfL+MhXwELdEk12ckjbzKElzHGSWzBMzswwqelM95r2g4uwpnOqaVyi+IeLH07
J0Nku3Nk3an3E2wUhNVb3wg24AZf+9kloZ23/QA5mJP/jyjItpoRK+dnqfs7Il6VH23Yu4XC+MEp
Ug4TcqjTrE0T2fEP7jXqJu577hQVeudRdISyB9jb7dMs2UO1W5eaeKN9Jdc2nRQt/dvPx2Ae/Seu
+60ey4RMFOOLlo0Od32AJs6QpRwzNBafijDQJpDepQb6LsLy0Pgh8pY9tfySQROtUO3xDyMywaV/
LhYQE5U/KsxbticBL3TWO91fce1p+ccnhpkM40fAzBsVYAiNxU6IcUngQPhuNq9DgpER2khC/gl6
PeZQC6k7X3I9veJW9cICwJI7nlbiiWlyng1tLCTiflEta+cBRDcRObARIRhCGFJUc29w0PjIb00z
5T+isJ3FA5U14SAXon2hdP+DU9402RutVqPTKDuZdSL84HUrj9KZw79y1w7bsMeo9FQ14kNVfiQS
W2Ow6vmSZRMxkYw0qGK9KbP/SsH1JL7e8IikIQJG7Nyc2ZHT9lwsMeICEgPfxFRwqcj+yefZUB3R
3jl8vu61CSpjcH20aTLVNPqlLPMpQtxov6bZUEJey5Z9GxhurzWC+19iE/7hVe5bPah94p54Q/Uw
DZI7SYV5ke6xsEG1vYaockpQCEgg3gXTrusdtKyOmYaY+aghiBbAxlBzGQixOfwaXIzyChEkf+ZY
DRTvUZBduDzXPJKOpd2Cf/Wf24jn6eAvF/G4AUqYR7WuvNxm6o3iwEP4xCofUSVygc26pXRj72j0
1HuCWbbRs9Mt8y/UYZZ1f3HWiDbV05cckfyuBIz7N5vnJf2e29TBOSrtqA97eFOBy7EFGKMABR5D
nVwLyNckAXLqBs5I7fbmIWHPi7AavhKp+k73vd2UsFtKzviY6/783znTkVwZwaJiOcfIz1Pp6UEy
jSuOuG0uq0RUtvAgBq9st2bdGCoO98FAsRXQp3gD9aOR4wS3XurT7DMW2hbM235Qn7Fo0dWn+SyC
slqhrUvrBjHyYDOE2T2qblqM/1PVJwo4OLibgjv9sUj3x0JpXLhwKVDtJP1SY5e1aTqkTASjOwA0
i9/u55hGVGyuaGbGidq2s6RMz5pyLzIzg/UbDmQbcnfGE2GRy5a3ALiyQsYsEeEf3jE9+t5oQk8e
Rbik3Bp7pDwMvs2UYW2TOU8Q0BH++/u/RR+p1/EwCTGbYm8CokbzkWsh/oQjvJ09aiPxgS6zN2XS
U2qxif7N29Z+OrmCUEOhI8GJ/cHrPMc9KDJjUZlYBZj2/CnCozbzurX27Me4c4nbW1AwQMNlv0/x
8LEiBQRgTtjeEUOuab9aBC09ze3ikb+X2jQtBHKLZcNabSIUZZol0C82R83JX9kGJhRFvkhPCpnQ
w9lG6V2Y8etNYq1jxbCnz87xXa8Gzcw571uFUUDrv3V3O25/2hzyi5Y1A96RbH26oOuCZGQWa8Kv
D4jwCtYMouuYzhBqmQ2DB8jRbnJuC1Eit8b2iX2/94VomB/yX/Gb6OEuww5tyUkzCULxobuAEUDL
qUQkug8urS/1s4I7+ZabjKyuHvJiNeGwALAwKhCpzSugvF8CAtm7AdFR68VSYEcCvDtVfn4tg2QB
Vx0xqpHR0z80y7HYqvBGqttVVJLJI6GhOsLjvi3otS2tvU3kLhPI/2Xws2DHlsym5ipXUvh41MuT
c9cvmqVNZ9E64bcsEzWQ0ctYmApv6JPN1lASOvxVV3CRzCd0O8MTK0ki4Z+zTVXLehyUOdMKVao9
LQZafVtcCrJ8SbfTMvFsidiAS7J32EgDYIkRn+7CLx5ayV4r2ntcZOFmTD1Dci2VowWu/FjWugCO
6uFsLtUmC7wAF5mCoDXQvpXoURzBKPwCCZJ/P2kbRDN860r3QhOShrPpC1h+WoCvBS870Wu4uENu
JY3NKDgUkQDpwCEmIMgWVRldXxPKYS17O6Y/mOGWDILi92nxdoItSSLMgX7Ee5pV7lLlGhH9sRsv
fpExajsviqo7gSNwLykcGFqbfeKm3h9cYQzSd0QGW+dOyMYb1J89RcURsAEjY8A0w4CXsmufIwYf
8F715FVPn0RQ1S1NhBXzRZYjU/yNsOws+nu0m2Og+5XsycQGPgeeMHZ+tqiFjn1CIcnm4x66MAYr
rh21SPvc0TIOtdb4mcCVzm8hcnzLgq5KF/5l3xpAQV7ABrSy93kzYPJKZGtEb/sLZMp1PoqIISDm
67SiAs06GLBcTGa6AWW/SLwEkWz9SsE9Zi7Dle44Z4j2DP6GBs52379wzO6Dr6isMrTLwd6+Jzd7
gZu5ThIMqQy+op3arca8T5MwL0HSQW3N85wUUnt8kz4K5Rz2cWYL2/i3e/B5vgKnbzRmd/qzJjx0
a6kKg37pDQxs5DZh5JnYfu17dMoZBrhh/rISllWeeX9TJ7swO2HLUY4MACzhzM7DY3AY1tQTHwH6
NaGYsaH27WPGYZbD1PO1n1rruEe5YnF25psYMrd3cb7cUqZ1d9oa0VGJt8NEjVZ6jAp3DxCFYi08
3NXysBSkgVB0Vm5Yxf/JcqXM3GCb8UdDTg/FngxziP2HaetEt+vdqcqntyRaYuHJmOPeGYZ+D2km
GunsKBiqm/U50rXLmjSkMMhZ1Sr6imxBghhPc1yb7L42w+w45XRYWbhcRaMzdaj7i0PwOhYP04Vc
jLD/K8CNohNn/LWs4TnB5Gq6QUEf79yd/0dBKvZ4r6XvxwjMIXwpPK4uzrGauOe9q199dDKLHe1o
yvQNyR6ljpIQkdyCNcWOrooeh2lhj5krNPqeplnjvT6skHYwVNF7ZCZuAw6mN5daYP+r9AUOBHe3
vFy5YZq8/B7lP3R//AVLFQFJCgbKgyqv+u+yfzc7rKxGhWFFuTD0jTLz6R262zz4Et/QOzWKjmB1
G3THvLxzdEm19YT5Yo8oOGx255Sg3MnUzISHDYzBGFmYu2rF95AWUMnBGramth+Z6UankAK8wXUb
0vw/P8bwcPdd9AZJ5EiOPPA0DZVvgWZIrwYPEKlptPbLAHYoFxj6snwqM+xCkoqZIE1BXKLG8TJF
hcMfKG+6kKntC/qGrcjJUuWA3UvbI2O1Q8mvf2U6AdZvh8ckuKdt+U/8PvLgATEg6t2gRKg5uHvp
MOWFy1RSyG5ckZ7jwG/31jrFOuynZltinkK9KCq8UQeaD0ErefiBufOJ4qsGM5k4ctC0mtA/7JxU
RsvYF7L/NzmVUvnLGysjkf1O/yWhqGwimT2VYH7ku+vJnNzutWct+/xAItQaCrrcm7MBLCr/HBxo
Z5s6Aq3fPyNPGmqlKAfagDHYFIeUTqgJ5LZ7g0HBQYRMfMPaJ5AOLZ/uRTPVg+Ke6m2DObYbwUNF
tW6Q5v8Rftf5OuJflBwz6YCdCFR3PeoTnHQTdtZKxg6NIUsY6bIv1Uxh/cEUvuRRk8NA/zL1tjNY
3VXEDcEnif4691cDuFzs6XNHwq9nS5y+ighraYYBR73jOPwglLfvWzx0OyBAfva1uQtzrMFec7dg
eY6DATJZu/NCE0Snbh7WXDU+4+EprXvPz7ycUP9hzJ3h6OZ4ufC5ajUHL7nR16jY6arPcY+e7Kas
M7kTLwIP3OQxsrjhJcFdXpx2ctbabK8ZaBjyUyQoxeu/rl5EvmDl8trZClHdpTUcXN4zxt3iXhC7
IsjSJrJtKiWm+cLX3uIBx3vXBIuDpjqY0/2Ey2AcYZXkIzcYS1RzvG2pC4ihDIsmLE07BosPBqTY
JYeLSUdCyAIHPNmYkX+plLyA1Pss99i+6bkn+f5LUX3uSwKFE1+TUAzfgd5rEACkAtI+ziAO3oMl
xU6xiOMbEnZfZMAjrAHnVlCTDColecoz7kWi2wYxROmeA9C/kjMDDxoECt61gIpxRGKZ75Mgs3d8
BfaK5hoSw5NtzSXfRS70+SwLZTj2vqa74Lc/pdJnX8lduFmDG3Oh4BCfxm3/guYEjcYn51oLQCXO
YG9O9bZ+auQdQVxiIdHu+LfCi6VlGROJt5E88oEgGPN7bgqVroH0o2JLVUFKt+DVpx2omY6DK8eu
ZoC8hNg+VRRNGB9CzofNCLAYESvUWgV9nMQuhyefFNlJurIofUynLqeBGiLjqZouSsar/O/Dh11U
RrSqAH8fqrU9lJ+ssjRFVfsgt+o14KDr2dxUkkgrb4h3YqXRYmDAbtHJC7vTvFp1aNYEk6yfxky9
IgBNevSRcFJP1RPXl/Uo//9Vmu2eRsEQyktGBFzwGO4bFOciaf54g9lMbbYDheToxy9XXGY1j/+i
tyxzUGJUn24shQlovfQYr6Tsj7ZBVa4zEVd5iNdkZbwy8uReybPKUMZLnioOZUEo0+vuhgXqCGyV
y3/WYpa1hGdtHrvm1doIN6GHEMedWIlaWPdZ3vgh8/HZT9EI/i2LySGkVejItwqWbwkL9dI711dc
VspYgNEPnOXz0Bv/NKfYNinaf7NoavxEpEDtwrljtl2/K9UIfNTAVgvEQphzq9w1NkVzqlA7DUZd
Xp6Uk+wDHmS7RVR4aWvcCzKWSeSkKr4r4ZsotJqMAEEaumBSss60IkE0GBiE9L9ZZ6LKlfm47Yz5
DHf0AZbmJWFSpzejqFjsRYQO7Sf4dNFjWW7PzdJ/dG7UVz6kHCNGUqgYM9M1iY3wdC6ib8mY7frX
sUGOd+OfqpOnFgl9DiW8WWsBC67LejE5xkcS/J8dZmRc5+qCw2HesUIv370vr0s0FGlz2JLrRlVd
iF6p/VzLpSGcY25oQyCY0fDX4z9qHU1Oy9bcwuZDSdxOR7pMUJ2j3orKzAfBzyycxP1lzSRRHUPN
w5v8Cp+fEk8hjqIK/FqYet8TnH/yV5WzsPK+Fxo/S1WqI/mRdnFRA8bAKW8haEE5/ZkgcI3Lm7Ft
+8tYGNTXjcmBDzyuaucQ82MfWFlW2D3Cs2U6GC9/oHE5iLzLfQmcpPstdsaG6DGnGXKgaMS69AHi
/KC0ZoQfkLqDv5OHcBzywmtx0hRo1rq9MHG8DqxIukscDZWCfS2GYjs0Lm6aXYCLeMNYwQVpdNSw
g+gU8KC2KxLMyF3cOQN09BE4LH2MGILJujb3meh4PlWbM/Tnin/dBOGrS4muWRxpTsL0PxN9DppQ
TqPGWEsm8OT/Hz1PXVFHNHNOZsf/DzVoGSKFv4YKHsYkqtPa8tC6jGjdbUJFq8C+FxpGVvNsVEs4
/rupOkmM4LXKIV34A6DXhF/ND8ECwpIlrWuQBHixmXe2f4cyJOFIhHn5v5e3sAj62YODBe1ACAUX
Y1dtRRqcyke8z6NNJ+i51lR4OJx/erv2M9VYD8wKJWQ3M8pAk1N+sqGmqrX6Rjk+ek/HcKGs2g1E
wdDL+DsjZdkmsaTgfxHmdS39z+INhEEYZZKMlFrdsrpnfrTuFK2Lkt7v2iAu6mQLz/o8qp+Fi+gU
wHCYTSVoufMCYf6X9JgDA0zYA/VS9AEBDaUYydWRdmkNhNRAUA/sUfnS6uXSctyukTkJaATDXexS
FOfZC4aSDOWuLHpeMWb+ORrcpiEYH+2A7G6J5DNjpL/SZFlGplyOvyeZ3kPD+blZ++8oaI24O3Xp
QZf1hJQ7yY31RSzw64x3EGsu5F+Uiz5amgiJ+DURRdpMuBXvfJUFuAakxdJ0vdf76zTzert616m2
EBU2etWpL3NajiUc4cuKBsZllkAnGO3+21NWoWn+1eziIwPuzLjmOgY7hTJg6/Ds9B+V7yi3aO/v
/UFdbCJEvuakg6Hsam0V0a9m7Vq6JjywMQGQecdXmHCKBUzaQe0xdO5mt8VJoLWD7ZOxvv85nyBf
Ku6q8EiHYLiDRiXoMKYUkae8yUS8VVdtQmIAFnUsX65695zsmxZ1NWJQNE75BUR/dqB5ip6TBuuU
9MXfCLMhOPoBpcAhXlFFENapSToM/fyLyXYqO6doZZFNBMgn1yDxY/WCAfcGSs8h1Cil1M5McqB3
VQ9f1XpUTEtrBNuQx3SH1mzMbIOjmajz5MjieQSDwIAkhjh3DiTDoTq+5qBJ6RVHHHnu4loiEneb
Ds6KZxqpJt6VA06KDpn66gXC7F4MZkarDzDMdgJVNlIHFA4rfTKF6cL3ayXiWrnpIiLYP/W3sGW1
Dsg40uHwINQq5FC2aDLbUq2aLikkX1bUmfQyRmFrDYth0cb+PY+j6RCrGbOWbWookcrW1N5ipZyB
9xElTMHd4v9ehUMvxtaLDCRHsVMjHXLbWZw/TarFhkYoi20074XkxK9tdyTkYF8PEKZ2qJcrQMS3
K3snWRb2xvvZwmqhy1VZ7wgXHSdY/7SRk2bs0exN6lj1Q9gAZ0co50ee0G3M/SRRLihs7xjLVg4t
gLOeaXq5d8YsjcbyPvKUr4c1EC/YGAKFr+UHaFp7fSEg4+hXMhSTBx0QpwlW84b0Xr+t8bU+u25f
vHEpB21PPqFclhH2/HwCOIP9Ncajw0KaW38Ibd83F+PV8WuIPkDuq5ssKPajjgoE0K9S9FbwqEqt
VZfXCq9L5LabnTNwhN7NpKGNYg5OfsM6cnIc14JUVg5QFaU7NAl/of4uH9hRmfrJR91JIaG9gLOy
W+CDLYp2iSnwRGMn6RFwTgsSark+saD9XBunOEvNSDicEDiLFUAa8pE8JhVFPzccn5XKVGdYzKE3
kQfvQYnP4zwPMIBy7aff6zhtnIEz8E+e39Z7+9HsumSoa0keG5fzqoGbSAcWkK0clfan05GwY/bf
yG0dAR3on5H9lQZ0WLzeiCgRciHeOJL/MnmcIk5ty6kmMa+t+zEz38ZiHuf8VTTACQ5SjFQv32AX
0zG8Axi3CphRgjeB1ws2cH/HW9x4vMJr19hWD8dHY+6/nZb9pNR1BFQxDDW7VbmszzwbCUAl6nNw
rMJhvnJXnKvfpKUPbaHWHeGd1UtkCVQtEpiO+5lIFAQg1YFuw21tl5sY1CChXNbOTewv1D/x1r9f
Z4exThNQuy3w8h/i9U7n2RKX5+ZxQX473jvjqIDVf6ZdT5y5zq53ohdKMgjWphZSyfJgQM3OCn4z
TUh6kpe5tUom+56bXkujEAhHD3WU5uCYP7DH6MwFw+dbDdZKV6tIyOXDTg7gOD60OO4pBs7GGshH
hH/WdA80Nh5KXeWOHZVA9kcJADthHyIfPMF8DXZ0jnieVu8ne6FTY6Res8HjFSWl3oDnrIYhtAPU
Ru4FKb2hRAXw9/F/7VrLX8HhMVC9nRqPwfaHX+zVtpCgrYUTQPfBXH07VbgihpEJ+GtFv2TVH0V9
OE5ifq8mYfFQ1RjmW++gHjKl2gaHXXOhPqU4DtNMggMORFYJ4YUfZaDVpyMnpIm+NWOkvmpcqytG
4SgWD/couCzgDns9kOn42LErMAp3fK6b2HJ2aNfQZuZtAKYlqxtcAuGHf+ZZ4x6Cp2nhtjR2VSWu
00mRwUa+b/5exY9N3s0wcuQQdQlGUO6s2Nlw0NkJ1sHUkPByKG4SBDGqSo2mYzuio1BMKEVjwAjG
HByfyOfc5Jn9P9ADNSMdxu0WdqULoys6+KTMU+lnvi9rBUjozeD1mPH2obtGWh1Ea8zEf9SwUYaW
0QF5WWMXarAe/7XbTuAyHlOkeCoHBaAI5SL1R3psPPGB9HjrGZDKKryXG5HbokP2/DsjYfoeKn9l
nAAsfcW+oQW7Sur2XUJnWbfePAQul/U4soiY7b/vHSubu7m+lYK4bjy7KeBsZRX2i/To52jVtaUc
zchyfgSRRrZGGVQ2kZDJT6+AdZ6WgZOTZDDd8bCuMsMoIOWs08oFbsyHvIFHdP5ctimvwB4sANRE
4MfDDBQ89+oX3+okzwoxRaQEd1LuWoDp98p74dT0F43UfZaGVcenJH05rKnNHx4rG+vkceS2kmkj
AK3l37aFQG7s8EeMPwc/RWBQjoggdRKyDWl1oeik0F83WmdBB3WlKHK75DdOoWsL5N1FHuWEbEGm
N6PObHI6OFoXN8g3qxYRavnPbbDyRTAZ3XgvwBJ3EDrthWoO/i5o8mFbNAKLHkUk+SiVNPhrQXgb
0pc3u3Q3g9kWrWA10vFWzLj5Wh0o6IK4q1T1UQ2F20F7RlL+pYT3IPFN2Z66bFXVRhbTG599MzFH
7lxjxVOscoKGCjVF48qEAWrYhnBNRs66eIG31T+3yFjt/x5YgNO5W5dmpmvtOPoWHyuf3+adTX0I
op95fAwl6rgTHgdIFLxHfTLEJbND1SHO0+204fP1X2dS/weqjizXGXMLX8wXu0bdQbBXgqV02SFK
X4BhUX98NRote3DncCzaO9V7D59u/njO1B83YpWUHKWuE4lEQ2Hroj1o0ceVfeZK9JtrgLABhPAd
zf0ZpbkrWbwrrbXh5i8eyH+/chgeHUCXYJWDhVqIF2w7JSN8OS9NCfGpMJh4IUIqMtNSL/pQEr8S
Ng0+GGi2sn7zsjQ0OtodNbKMZPCYAg0Ro+YWD3z+K1hDD8At9ctOabN3ctBnxm1Aak3RCr4WuufG
7hXv97TreVjDoKpImLFzsQOcgPfbhRinARm0hUELMdJZoXhq/3B3r2WfnPsX21Wky7QTpAMo/2+5
WLYxCwZQ11NMmK559kR1WsFpjdXK/MdggAAT8hQ9TZvn5EqGVOEx/NXRK1OmiF/vf36/t7FQzP1l
oA8A+TfGYCui7xli9Q23oKnXLuhNT5LHjH/b9eXXYuxBJ38ONn3cMGH0JH8lyYwTHCgQa/+qJxS4
T4gvIc3Z5LVrgM1melNa/P5C/UcxaK7gqkhhJ4qjNoNhr2owZ8Q1B+7Nk7qncH18jMI4kT6kwiU4
7FZrItHVO8/9Gskp0qNn6NMf50ube7j6WVyVr8jci4XRZo3duEU1pI0HBA3WxGPmZmXadQ+Mcm3o
hztPg2SeC4kdYKhIm1NTebu0lQBq+NLW1CJJApo7b5LUydZHCbOe+kG+10fUaD9ehegVgooLIxCc
Y3OUlpkb/tVd7v8wf1KHmTArLwi+iuJhRvKlALIQSjhbzTvk+h55+AHijhys8gU65+mocqseWydZ
C5fvZ8hRjbPsceS7l1TMJXSkJpgW0VeEFCpMhBkgD+hkxn9qfQy+Y8uuL+8Dxu+kS/sA3DLyudvb
h2JnxxTN0kB4HnAnwVpy1I4qQq9cTeX22xZrtEsyizCf09dhcxDmzcHo3QPimL/yYNhOGR46mnI7
ueYyxJ/4Z2jWMUJhWe4s1X8FStvYrq6Blci94N/0NJZUqdT1WwvuYeUFwda5Q52wepEZIzCqHvGz
Vas/dgubB9YkNcR4c42f+55KmMJ45fY2uqR65hXpfoW3jm5IraGuCG9Dxn1bFAVbkEVHLiIJ45o1
zzFALDIacbqyhIZA/jFAjmJpZ0eD77wd9x/3saQkGJ1OcwxdDp3HWjjhr1w4QgOU0be/cvZwF1m1
MmywwdYMF67hkzEeDB5ZNZ1i0fw9gMtNnG0C+/TjSFr/gV9TiifvW3CIFCj9kpgq3vY7Rr6PPSYl
v3+eaf31/WYJQ9jBmoRWegacrnU1yxs8tq5McY4fD03lGe2wqsMLbvp5Tf5N3Z6WOuSSWK/fKmug
CoYRR2hZO97BDHqQHzg0NhjpUtyUgDSKkR+ZxqfFsdbP+sOFkAF98eZPGsPHS8g8UOja6XQfCNJe
9/YLkuEI3O3RrneUcSaFuBMvJMaHwPBfbWlQLyMTINy6jjHh103SgxHf2d20n793cRAQa3hsi/h5
JZgKdHa4HPHV+ZA5HTqE4yrFj0rEf6Zg7hncheWanVq5h1WDssreKZzurRNf2G8zdHcPogjT8tEz
A7HbZb4GxMInbRq8mLRhtlKV7yot76jq5sl83GXx57eckWnmYlaIxVJEzYnR9SXTENIpgdRuvRN8
MDD5bn1K6zTaedGSFSKrLIZq19CeyT4DEZ7jtc7v0iicMZrUYQvI26J33oRE4dFLHKVzkGyZ2Gy8
Fu4DRGB5iwH+mjHkk9YZQtk368q/nPVWKzoT/nUOTePgtLCvPdisk24wl795Fx1rAPhD3m1u2X0u
ZtXsdNyRQEO+cuXAcw3nsmMdtF0ab66jpXqhnF/KaRqyhXkDFfJhZiMuxJ7/u7ZnqI1a7/5NccaW
eqwdooKMCwofVYyjHahtJGJggWhMw6D9lO+QjqpSkutEN0XR42oQ15Nuj5MR+pDNdA2CTQxu0uYY
gIzESyCeYMZVYuTq/wnwGmUnx4VOucSYy3ljzxUnq4lm27P3DIO3bfFKLioneJBMcseoFytW0tdo
JTRDMn+7zXKjObEl05TwRfCigcABd2OKWWvHVB4Jvdy3CZmQozfuRMMHbjLxalJTmhMGeSiRAT76
XBi+b8Xytk8PTvk8Olsyku7+BqnnxTRvIM8NtfesIeir0FHC720dzAjexgSgOnMub++OFj05rGAC
xseY4GwCH7aIWRHL/bRW0Sz2mKxYqPTFeQcaMPcTedYuGgbdIfCyoQB2hedFhqiy3OPLszTKXenW
5ngBaHqZ8nl9PxAi8i2K3uHH+UKAn9vQ90QZExJt8txjJ60a3sSNYHof5Hclz3guSZtWo4XfQjW9
IB+ZCtFPZSY9oTcnoPlVoqPFNISZK+eox8eYzvS3DzFDa5dhjkvAJVzYHgjtrTR7nmR04jAs62uZ
wViXiPPLgFSMC6RsW4uEaoe45cTTRVNBL0KRsPKnIOyQfwYQC3ei/mZF/k4M/lCv5KzPIWS5PaqK
KcmEwnl+/P03acI4+47BUJMgoOGm7eRXONbfF8t4Z6P8m2+CUXYKmPzmtEwjqtEQSq4sAbJ/WVZX
/F28VubPRzECXlB4HUDo2ll7hUHogYbv8pwEZSaf827ppB7ASBUnQAj/t33JPRplC6ijSDj9m/F6
jnQ5TQ71IxkVK+0nCu1QOsVF2pfSQWchllSMbEYQx7ZpYTyn+DkF9LVzmR3LEZA5pUMDHyK1kvhT
9J4WswuuUdYzjbD7aIj3OPYYGXRUBbVi6dL8ypgkHglFVBQefYj8wCeEFZ24kpQSoQ11mGuC7aQ6
f2ImuEQzY8KUuwjIynQqsGL5OJC6HW3gZmgSe21h4286+yO/g2KpYElsK/eXm8V965EQeNZlJ7wV
JM5VypIKJw6LBIBpLSsJsYn2CbkVMBMN1ipMQWlyZz7PMYUe1qPU9UlvHN0Lz3PFz0wRu167nQxA
bSvaHPcEZuoQGTaBnzCb0hD6C4G0Pf4qF1SOFNNs6dHaoq53FECEnUuZdHpGWDurPwT3RqQa6moh
7hmOixD5gkly8eGrbtLn3VVNDqtSvM60yt2qxFJcvtGBG5wNIaLfYjjhannxvQrPmMBZDQ+YVA79
W9YSRiS8Lbt31AWdXwdnZ9j3R/MVbzG3aV/U4IG1nPwlj2JF8Gr7UKsJYY0xRoRQOvpqYhimumQf
ZN5ZsJOqrZjv57WDNTzJtLs81etRz5ZnHc+qr9W0CJyVSYzqDV9ZjHM42Vne55ICTCNfeo8RN3bW
v0jR5J6hGSCHx8OF1XCcLfYoHBq37oSlJNPCmRcX+UEVJJXTcQajUFAmgKjO/3ZpNYaroE8nxI0L
znaFGWCWgApNN5Oe52f8Pb7lokio/iQCtVVJuySXfyYaQ7GZZLpA7WoFFinoVym2t2PFHqDRO1er
yQupR2El+M2Ndz9f8shQQy1Rb0bQ/XG3N1y20w0R4jybQ9B/TFr3m+x287eJ1q9biMgjqcRm51Jy
F1yOXrktSNHcAWq1ZUhEkB1+2Bap3OPRDi5HJbgs1ahb81uxGgllM751FB/5k6ZDsNbZS6DkrJYO
zkxqjtyfmiSxSKQhtfoYI6i/n+zi+/j8VEWt9mIbpAXspz4VvWRomTU5PVyTfZl1+3IYdjX6ix3S
kn6TFRbaq/ltnSmTjmALH/tUjwPvJRw9DJO0/RD3D5VUt5nFHpTRRD3MMEl2AFfHz7LYe07ClNZv
0THf6uPCIcvbKn+EnHlT1J2svoxEyjIOy0HA3+nDGasXConmUu0lVFlRSNjb3zntoHjXSZ/i9BdN
Z9yBNNbxBFb1vuC03Hmv0Es3egK3/4A+DC/v/PdTRJ5nYpBu6J2YzHYGl0R4ANOE5qQawh/A8ImL
VdF8hlLGXPhFNsWHPeN7Qw12tvT2uSnM8T7VQVTnZxCztO3CsH5Icew/33Cz93iHIbU7HxWDJpds
U03wsNg0IYJJd3cDJNIqMcqWm7IBtI+VxlVTpPn2x6Cx5Wafu44Kxqqd9nMbe40RsPkB7uqPvFHr
0k01eoHZKfe3q4dW0cSMgVfsdG7JfkGVcfNPU2pw35Uz0q1wiQwgu0NDxmF4bSt9KIyx32KfMG++
GAX6stHsqrNiCtLLlxzD7bDqfWnF1C1o0saaPlzo/I16vH2CXtB5yYtTnOs4ZYCTMbWq7F6zTCT3
nALO9wkoazNZpgejzTFTyrAoltq+28DolWspe3Mqj3t9/pJPj7wkbTB6Lgytb1bliuikovJGSoBV
/ZwIKOtb2Cgjs8lns7ld5cGPRPROyFRGN+mxumImU+0/JbcrmQSqZwdmGKE/xvKh9I0OmvT+0QTh
pki5rChRyGLswFU2psprFP+aKCHE/+VVhnrQekDFAGeBC8+R+dg4ynZJkbP1+2Or4FPwhE+9ZynF
0+dKYgFK8O7da7/SrF3BhxcggXW1DEaKb4f2xqojm9dfUrGTHxr4voX49HBnypQrXMCrUeExJ3Kx
XvIc93G0NNSc3+FZafofIrbvoFlXjVO4qmuebVIwZHFHGzcPcEN6SIP+2TuCQeMymGH71uRdkiou
6qg4IJ934nMcir5j2SulOW+V9pbBw7hCfWU/Ww6qwCHaQ1cfB3bJahUxWUaKRpO2TKPkgEYlTwiY
9lTI87tvLNgcYHHmWK7oTHrVrz/PNftqgPk98UYW15tZ7neGoE1scCuAEyNDP9/M8w5oU/D7XUF5
AffK9xQ672DSRG5uf3Rp/fjRj+9HvnQmWniXXz/2iV97q/hnQs7g54B4cT7wn6u4uaqgoU55bkvf
DHCurXee9WLqOoTWxEpsjYOWDivMndM4sS16F7WMmQGrS4gXki+ZcYHHjrSUgwbb7/EnArbdcCys
YcK2YP9SIEg4esETRAHFpYyyu/zI7ARKacasik6TZCaHBWYfJNlzvMexUKHIdvC+S5AMBNYKGT2f
M/RrcrGst/TQJG84eZe4Lq3yVmDgaeU8yDqdWTIuHgajcHRoCtehk5EkxU9Pr1nJldmzQ2e6CEwB
wCB2/F6etzhOgJbwNSYQYBjn0DgrsjhGA0pJwBtcQ+gQBS9UZgxocC8RdOzWbZq3mTfr5ZWI6rcn
GFUfnvo4dwhiRSyFJV6nnwOL1aYcwOWz9MkXzw/Zifm7TuHmATb2JhivanTpUF3XIAYr1jKIC7CA
ZUGETR6jYUCp0ZVDOSpV+o5ZxBpgMfvAbdqihFWMoicKJY5Ji9+Cy55ESrHx0x0prcd8tvK7VWSx
0i1I8sokXqYQGruYtgqBpK4xYITo3oDbp7Cp20qADXgowUWTfiO8DhkjkUfw9FRriV12AxzJxLJe
aFaQiiN8e5ZqSXQlYtyrD7VlhUNvf0xRvauN+7j4Y3wDvne0hf1+1zTJ9eIok6K5cUxHWu3QG2ES
kaVo5iBuGnpwiUaa2XfIfaaihK4I609APRgX2D721P9hTP5gXmwSs1Fn4lLQtwc0OT8x2lAqr0L9
uB7Vp2Un3uC12Jd3lX1bU5sxDp3trEhJLZatm7Ln2LLEsUUg6P341NFKdjAzflnYnp54So0vuy3Y
lGWOYEsCYrWjlEc2ttqpuYopryvLscP9Pg3Aw8nCEhAICa7ZKw7Szll+Kg5MWHKdkX4VLQRLSPix
NI5dFnS+Ujx/bYN1eOsoLj+Gx8bCf9wDBsdKZ4YH10vA0lRu+jYHU/dJwbBlBEEEfJpcGf5p+b5A
Ov4ArnSkXINkkfdSYvBVnKq4fa5HNs77p5ChGhaMK5xn98u1LY4fA2i+ytqxMHGsOoiSUL+xDWLn
ZzfQH80DvvjZA9v4wHkXVOSMg6Tr07QyZRt4Kk26AxfO6M/p5lrAzcbJ66sgGfH62IbHt3sRiU1i
oFvpb9Pnj2g6kpbu1XmCiuFgq8Nm0d52wY+rXEoraixBaezTW2c+7f1V4AW9kXXnOR2ri5i0tpHa
05WOcRWXh73HtMNQehAJ48MY8voWMw+p1EFhaYXAYDK1Liw9SO4HE6VPwOXX/1ACqpXHQ8tR7vsR
QNhZNgx4D/3JfoDMbQypLKg+GBtHvpoCyCGiGU8TKbJgZt1XrKECezL7hNq1TX8qiEHBe0xmyf93
3zJkBniYr2i4lYuTIkUNq6ciDFJfd6Y8Pikw9bTrPO5dzRzHb8x2/oDe0vhiPwPXOtFM+06+4bTN
jUcwgu5zGBE/kWsrgmArOzV3XUacUtk7mKjRFAAjnEnRQK6Qc1IXxooeE8cs2i/okvEwDR8sh2kU
OE5pwluae6aehuHFCI/J3vTQh2prUWYlZGphrABoBNtG4v6NeA3mqUTYCgA9fh3rU4EJyd7E+/tR
dW3RvKAT5SWXamcAk3RAI/e2/sDu2J/cLR38eKbFGYhrpk6nYP4ChECT5iJ7NN5B23iWb+JMVq3y
UlF3pszjTO66ZCyqwKZo1ImW+iahoPEQQi1VKZytyep0ERbe1Slu3ZzL1XZxGY5iuFLPHXOq7SXa
/MBZ6fgyX6yQVqz9lo1QyzpQhk35vF3DpgNfuS0+PNeTKWl1zTFEZYtXHNc0YXh8pIl29mH6D+RN
WfcB0oLsCGgwwhYU/UCTQwOaZLMYwm/5UD6rgYrfbdbeDXEiyot2zATrCiw28Es4UL1QmKCw9uqq
F1KpFGMNKQnN+QZqbQjNgyyJzeB348r8Q3yLra47xEOE1jCUGh6DrWwe84Ovwc998ctiIkKCeSq0
hehG6BoQJ4kcQIldM5lCtiS4M12MwM0sf0l8oMkkyr6YeOUDHIRFkd7YK0DvXlExPiftFF7NzPgJ
Pb8yCqJ5g02MUBwDKAus+724zaYSPdWzI5eByYIUciSQhll8CsMXNoYq3lRU05jg8eCkx471FS/a
oOfaWP8aGFpCdAcAoeDmmy2lnzs0PaMllPm+7GXZVgIZJ9JkvsaFT92v15EBJ859Cxgq/YKb08Yl
RvOd58137XP/J+OaFoWMRySYBY76i+de6jrX5G98MS3sglFk6w9ORy6OTrKceWE5jhel/yps636G
QhdviDeFhZBFk30ZDa3NZclbqaxaSmSGQE4o/vfNcnAkLUisxk+q5VP4k5ivOdfN7KanAP+/4nIh
Dwf6fcKdJssphUbkdE6zQMkI4GsJGVfDf+gM6AaHaA7iie11unGluWg05uiLfFfF0I/GJkp6qPEN
01e5fkr5X3aPskhdnZvtWX/cy+6yEo41QfYWYN2YnUnuz81iIvdicM00LnzVrkVuXVXOVYu9vbG1
Z9e1xls36hyByKewiwPSmes8xmn/iMdSsoz0h0OgL/wxGdU4I/P2QGyFOpIeTGOUMvV6vfw70dXc
cTVhP9aFgUyRkruDGSMAvQaCkgNXBlwP/JFhUzlanlHqUQwpejpwgNp9yUn3do1zj6x0t8hugx/H
Nowf8pRxxs9c5mj4M42XwF1Mo486ob2Q0ONLl2NptMYUcmH02g3nojZw5tnp5VE/5m7SMP+RnzXK
LjteDVQ5C1xTXM9B/jTYkweVUSrGrsUVTbi+RluT3Ghk6HiNKR1ixEeeXQtOtem6PgnGVtotUNW+
yQW5uTxT8TABsWxUf7RgZcvniEp3PeJTebZe1auui1eLOZxm6wa3/LQvNexEdQ8CA61RqaZH5Evj
FyXuJoFgH9PfZaxKxJXqxkg+4EzC3iJR9DZl6onX1XSByNf6S52eSVvx3oXR2GyOkTkvWwJZN9Xz
BCwMzNGJZlP+/x20rO+AcwMkBHQar8uMpfayib+W+UbjQ8081z7RxG+Mct91dzkV+lzbUO73Nb+l
mFjSPfUb/ZutF33Uee8HKu67MtfVqtHW+Ek851MzCFH1oWRPEbl69fSuxvCUFzkblRVt8stljwBk
hYeF3eVa4najE83b27vahXZIi4GJTEb74wjGCOZ/khqVizA0Sr9xJk/whnXl6v+bhMyEidgraKjK
ghHNfKgLLSfLL4Tolcq/4209wvUimNYSG3q3ZqN3wkcrpgd/5hjvv8a4nnc5MpUVfuoH4596bn6d
OwYROjwBj7z6FOqWSHNC69V+Auz45+hLC3OnyI0aZEsMqeS/Wt/LvDm0ATrKxnBipKt0zX3SHl2j
tAklYmVqHKB5lM1pXI5XVOw7ZLgi7i2jvCo9bU72+dlEoHNq8AxMIlc+qp+dIYkQ6T2LNNjOMBl4
v0QhZlL6Z7lkV4P6O9sXAUlsHha6d6cHXpL2HdSGR6AfFd39sQWnNhrcou5TfEsFgVu5zPMZL5la
TeNNx1Mp8zBKZgETLJeL2nu8lucIJV4lFrrKTWw6qbR40EGk+DJubE3zULFoRqwnBsZ9vfFXeVdX
Os2s58Knv0xwBHIS+lR5UaA09PTzVf0/o97zFFnFrBioj7Zo7nimRblCdmV0mHuWlNz6zcS/VwpG
pOYWuS7QFsR+GqYnsjVLqt0XDDEmeBvEaskDvo8Q5sQEF4JmnlfQnklnvcSeyF0qIdzTl3xBFPZ/
GcQuONsyn4OCuiDRex3ODJXSQ3M5wGgVOGrxYLAgbMfHrqKJFNj7DA5nNkWmI2aoh7xEDR+kWr+K
oVSnm+yZD1030t0MQv3RU1R/4Josi3l64V2RXFd5uIXkyiRDCdfOOtPDcarEW4SKeXRHxTB0XMOF
tWqShX0xSzXHf/P9/pS2krhFRChVtrztD4q3sjy2c1HR6nl8yBf4hEGSPf6ofoh6OByj6pBgQ6gx
NXgWjBetZBlwdBdwZU/nu58PuRs2NZc+oS0DWhpB69vduUJ6o5mJNzijjjNd8ibM/znY2ybQsn/U
+fUeBwRXj7/dNA7rQJw+i7NRG6OQhT+wPARftjor1hgAGXpyC3DwpkA4IPFL0oUMlBXUrBS1khBx
vlkGPRsJ89en7XS1owJfqFKbsWxbwz2xcAeBSO9qQdQymgLjmAjMg/GcTf91Gp03d90Uu8xCyumd
ab+HxdbNoNZgrDDrVaXeOcP5Z2aN+DMPodR9UUa9y71UL8oPPKEgJY43et4WYDnDmV3fhkGyHpqj
SgSJyfPXjo8twyU2NvXFSHD94vvk9ApCsSXBmg0+BfJ95o0gdR6IxGpx8NVpJRvdVl/Jn6fdQK3u
U0V3zWBC1DXW1wsvpYZvtd25Q16UwGwaUCwY/0wYbvYKc8+u2XTdvELM8uHyNH8587/z6Bb5DfQd
wQmPjMpPc/xXo5BgGzv3eyaOb3NzeMD0pyaBnpNNQ0oqRqduUPvFqmKp9iKWiPTi6PxjA0Z/dBfk
zF2Fgg0c4N6BUlC63FpzGfoNUXdDlljJn52YMc+/CQUVQRf9zjMgt87SCpZWb4ZpsMsCyYcKrNOj
ND1vrTT++FqhvGhvkFEuVaoAbjFHkZP4NkCxuuCORyg0ZBMuu09kY83tGOfhYTr7qEM5cwYBgB6l
esyBYiRkEQ3tqQc2zXxldy3J/vdRyVN6PYstcAHKYGt1NmMvJxFw7UZWBkrsgb/UrNd6wR32c3i6
VGo52jVDAos31mPIZttbkmT0bcw35yGH0qn4GsiI+nEzWXSyDIJZaW2h/Td+q/p6mjDWgKpVZ0Xo
ibMv1M4JNQG1B5vFjzP9EyVooQineWcpMzkgj8Cp+pUhvTSIhMRMHimxmZ9ax3Y+UmgU/yAI/Tvu
HnLIisHt4npW6b9DmFeM8+i8UbN5yAcUx6xYK35DebrTJcQr2x9YrAcbTe8VoZoqmPCLsDOgW7+L
U+7HTERSyaAVwSI0G1m+/pEP1yuBbMWjhEgiVZCU8eVtgnjOrixnTiPl8cbJ1Po65YDfIA/iISKE
lvpfNhpxXEXBRUULOxqIJl9NTmGF2usyI7zsLtZyumT2Uq51J1RjQAaqav1CNoSOgrj6O3f4/xU/
zUodeoXrz0YFnA6/mhjFd4mmeZuzsyg75StFRpBOj8T1SiNnO2kf2WD9jnD/U/M303J5JGzM52GS
2BwUV9NlDb7L1SQ5AmQgJfLYRkJvMcxSVS3gRnghNffcXwrpzx8qOqT26ofMvpqKf0FtQxNQPPw8
8yQhKfC4RQsxRIWIyhtmNcMKfo6inYa+zRGg8UToKdYpjrI1VHt8n0uctP6SNIYeMI/bRXg0dNrU
g9Zvx9Bw9/F+WMiyTZ60eYDfjKHd/9qUYHs55aya7Pu7ftFeKSpj2ysw3bEoth/1ohSj+wsPfYXn
nLtnIcJ0qqt3qmFUIeuR/bvxGiiUToDQTP2A8X36kgMw4F+r+P2/PzDgIPDei4r5NeUSk2xhy2+x
03B9au8DEQ83HH+PpJ8H4q4pOqb1CLXaE1qVRu4YJlS/RPk9VKDOOQe1zlF2fV3nb4WaMaVWd6GO
9psk7DyhIs2HFdVE9UIeLpwPepkWMtZdZsfWcHQUAN5M/seTA3jSc39UsKaOvp+tGiXMSAi2+ETA
0r3vCIHLhk/e575YJIkiJeLcNnnVgDTPgitN12NKD4XiEsBHYiuegZc/8lCbQa/AhyUzKme5iT7I
zmPFohpSGo3XzpxdJgK6ItYeSd5wz0Ot8cWH5zIV5GP53grsXpXhdf9Z4gFv7HD5c8bxMFKLIg9P
j1dmZ1KsujBLgnniwlihTFtexdpyZeL0lmN6AqOP6+xX4/v5YYBLaLshmGmmcWR59hofhS3zM1Aw
Nfz2LdDbcIiy+oeCzizKBZ969HR/5TXsYvnBGjxQnc6hsszIWLOoHkxqimIauTYtB+OjldzT3D/S
mBNOGdWm7Xc9i2yymKqC4UTHBu6K2N3/o8ob5Ab9KpnbVnVnlwXTjyhRR4erfdZjBN1r3QzSeV1E
Yc5d0yboLW2w31EZ1aYCcURgERSSPUIti6tQfBFzrwcr+PBxwPnaJYcPfLzG8n7q6VhgmQfc4ur9
/+0D9vNHahIuuu1JoYVWOVF0QgE/LeDW7cno60jbm5nEZJn/jogFDFV+m29jYWrZH/4H3CoQKdP3
MsmN7f1Mc5rUDvr1/0a2O3I/pqzFxBejY3lljIYE7UlGsVVPFSZQ63+PJMOCLyi6lysxm0nFssJa
zoRVBHcimaWZm2CyR8O7PU2e/PypWeIj2yj/wxgtZ34hn1JJQBfGVuJuwth8/6R4FVLLG3buMuwD
wm6NFB2Llq948zoGpM1+PCBgr9FRgy0kfOxT7zEQxL2NCBJVGCXLzFdON7R9R9L8p2WTU42QIamh
kTL/ZJYE94KXxWlfxlxXfVxrb8iEHFWnPsrRGZCkMnMrC1x+Xuk3fR2WekaqWzDZgkJHPS9wGmJ2
nRAKsCKXebS+f9VIUTVPQgJjSw+kCCTjE9DVtsUDpqoyOyviR1L2M3XX6INz1WmeNYCUdmviJERJ
rRIoDEx3+bp+xRdEmG4Yo9xIvGo8mnnXxlm7m5uGNtAu86g2R3QvCS2O45/OTZDJRdUIdzhrnhF2
0wBao4QZmrHUdD5iBb3D7yeSl0eY1fCdhzc1YBGRbxJ4xnV0IWIFADakDLE3OoA2eXF0ce41VpVw
prQaQ/CeXkMCsot5uB802fDLgjTWVPgXJQ0mqhhNENOeFC/HhqIw7kFboYVhZOLRoiDyk1CTzjIC
S20rZt7h8ugYCNsFzcPmR5iXrjh5jatIGK/4IO62J+japj1RZNepKCaeVbR0cerOfznOjEiXqwsd
ksjIx2Hh2Yuz8M1kt34ba8dkUuyiMRuqeIYUMwGDSLLq8dtGV8+6D/XUtjkYt0rfeaE9I2rwJdYv
kDrTy8XMakcq+03mUam1+ewNyDSkvhuTxeHZiZg9nmisUeC4K6u8d+J+DIv7VNvjOH/kz8FrBbon
iEdRVU4BTmFm6BQSJo+aIcKuT5CJdDqVMCyc6hUYZaRRkjcCOOa09QDFzpUEq1l4UPv90dsjoRXw
lh6iJhw0fV4ecmKbVuc8ecS9a95rGiR2Rpcdg3LZ2W98YqfGUUuC87nOGjWZAMmXaqgszgqJV2dr
24vVmVztjwPORpARuqMEsNkKFjjBGv+71eYT4oU0KCnK2JZ+kAnSsL2xcrvigmsl29FzqIFiPf3T
b1i4NBS4JD5Lp2fJieN8el16FWHr25kTfL8DT0FFgxDbie6k2FiY7VMO3dJ3h05LAZgktljW+UV7
fcwrjZtv/kjxkIa5WTTQeCAzctjYEvs3jcogcuLCT/7+EwKmSx/uw7OO3fqeQF5g+SSZ9IxeZmWN
odWL2VsDM/fYtsTqV4RY4V8sysjkGUDPGzAnicWie25JNWncfdnPIbZHGw23Qmn9MlUD+08t34LZ
1CBRBOTR0Lsz23Fqw/MalasRRHulwwKxtawzCxhuvVXcqjQecQdvKH2YtJY3hBPq5lr8BlDyeBcZ
M8lqmhCzr9WnQ3Yqsa2uP/Eioxxf5liShZQGlkICym6LblMA1dHpI+TtqP1ozG8Q0XZBZQr7jPVs
9q4cehqtsDNquo+0Pg7NdUXHvYa+026+aIER4rfnFu7F/nS+tg83aa0d2MyrT/wcHWDvkSuGSao7
TRBK4SyCqvwlC2a7fedEryKOyf4fm1kcjsVzX1ojFChXgKS1DZMg18xFNYKrv4Ml2/2Nh71LjToM
Qux5nRWsa8QDZQnrR2o5pLK4OC3Nt8iQ6XW8u7QHHEpcJ05hkT0Kakrp+QMWNnQHgxcI/0p5n0Oi
LhmGcS1JtRLNgojMveTh0v7oBioDCiqHA7MQmQvcIhN6juShtoaNe+hzQ2TP7F2LZYJp2G6kWEej
3yPvz3PI7M9cGvdBqSQx0Ef0H1pAQ6qyVejqjnnfsxy5IPgyuZNdWSoynbw9j6dVmYohDFLm8mTC
KG3CqdFajmV5QO0I3xFKVGS9FuqQKVpaT8g7O2EKGudBhVz8Zzy62mEAA18+kFWYxBXJQNYkRs+c
woPQj/RkvPAfVwJGYw4ANqRCX50tgZ/syU6GxGqwaWP+0pMBrfO69Dw5XRX0gmp0Y1C6mjQcYQ+g
VrBe51Hp+eZrdMCoHymeDD82b58EVOqhD/wMolIn7WfWYtLCYqhoAovosvHFoB4BjymfnGNW8pOi
48W6KrT3epzevrz4i+GVjR1X/Pu7j7oabf6B93DThTtcbjekKVR72W0DZuDrlSmNJI6J7FtrYqsX
5vgnBcfQ1p9HIOz6id+aXtA06/AWnIon6TJpb04cSinktfTkiEfDJeMBRVZ8DHgDG4zt571kyQMi
cSGizJgJ4tM9l8pUOsYzib1N7AD2TmQY28Tr76Z03c5QIJTUx1fLlDDRr+8pTPK1C+tH0MVcPd2b
xfe/BO9RR0U2+5TCGnq0Al9bORsiU1hbBqYLqra9CpCaRWLAFh++0SySkK6e1cAwSY6HRKD/EKzs
1fgeZp9LELbho0aElmTXjGqSE6pSEXcF829/m0DsT2pRObSi3YQ7ptG2Uw5MK1qfYrnCOLR8uRzH
STsSmvRcTfj0x1yL7o0LgjHwoIEMBvJKhaSz1tPMN3ndY0KFzgTrMS9fuyhOUrbRLEw5UtxMADM9
Ux+oQnvZqBq0xeATT10VShbwKVdV9kqANo3Onxb1hd+Tmscr3uLicwP9Iw0ZXZVCR/ayCnxloFV9
LRaYu6IrRLBRmbhsj9AwMAf8MqZO/uWgPqPEQsG83AvaOTugU9QpwVc7Lk+dbXkCci27r9irk5xG
9zJnVHsiYzmTwJAZZBLJw0dWv5+pAN9LoOvfEZlzUyqZXfhAdZv149SuKrhxxU4U6PkN+vHX7ff6
U93lyvoK3tu7MTMxHZIc0hAF4xcXW6eucgQe2bBvQHHKjreENTwvJ4cSgvsxSH4ViKQGMQWwdx7m
jOhsKzHswx9p/0G3m88cWcbnp8CF1t1gTAEqE5xMZrjc1kgK7Wny2AJ9d/UK+n5q9bDRZ2x75R3x
nyc/UAGAaFr1yxRwQiciqRYepnI6Hdn0NybHrzKIij1I0qTU/dhrnZERzHJIZTOKgcvytxrZjE6f
B5ByPh8envBErM7q5oqrrz1FTkJO1k1hRbO2uYbMpp14ldNlga88YnrnCsF0y5VgdyiWvphenfq8
BGP57DaXflx0ApVcLx2f4nZHzQGV9x3CUm8tWX5UKtHwh+Nf/3dCqCxgEGEOsJnw7aNPptdwxB5y
m+Iixane90SN9eh5kO/O1R2jbp/YVmCjCPtayjkaBagXly+QQpfjCr4irir1kpcCgDJij5z2GSTf
ti5LueiTJnYBduojtIMwIwURzsn8IIKMYXQ9iro37/fQZuICSGB/456C/ATKmuOrte8hWQZSY6aQ
4nhgRhfAfV/vLYpOhO7MLOOankY/9ofaCEqJY81IzlJhuSZWWw6Y0uBDuB1ixhclGqXZW6FjhRzi
s0gN6BYMrrwtvM9dj2gv0vxEAVIfWBr4R2QjJCwAIfxWL2SR+5LJdlAKvnskHhep+YufmIVq/xEP
P1emgo8aJNNPBqSK+ML9JFgSNgOw84eiesKZqne5n7WJqsi85SQs7llPg9uyjAkvVGzhdpDTQxDj
jnARK17WL6os4RYkM/yp3J5QTtih4CI7PmNQdlGFW58VPC+3ss9DbpAeKxqNGM2gm1teDuNT/3Ww
T8P1WNsF/tA6szF45jyg167Nf0FJdu1WikGv0Tl5W4rrHJiiIZJzmHnyuv8SNtu6Hi1VnBLIeKw3
9TK3O09iKySVGE0LfJGc4usrH2C4z2+Gues9y2bmD+Z254EbiYE+Q8sWLR30BzitfIlKbZvJXC+9
8dNP0pKjILBvxvuwu4t7PaNkgjrwNQLKigZlpuANHCtEjhgrwEkl9FcxXeAaMNZ97ImYQnJsY+jn
Gu2AtY+yZUCmiNo2GlwXgpfTXhpD/g8kAHWmh/ufUsVxyUOPs9tpduNALZR8tBb0Poi4bXvnYwj7
F+eQMJPvhrHCuLjl8W8+WQBQdhZS/q/nJGc7o8WwOl/HkCcYwZE6i4JH2BHA1iCKxR64T/mhdYxK
rUajfuU9oVg2bVs6hguZuaIjMFIe4vQarTrw+cy5EmBImVt78CbYCOB873Gl+LH+V6ChfwnUdnbA
zqtCmPFiqw93gXdsxOnRgNWcdixze1vZURvL0mhkAfb7kYQrpBiYBphIZq3Du2ng9vR26nMzq9vp
jMMfrAAzEOvqkZ45fDSuoo+Sv2VXJ7FhGXpAAWT5PHjRpWPvKa8hwMM34THY8E9/uesDK8Lwz58K
WGt1EvFq1wFCWv4pdtdX0oAwhAhT0hajEguwYIExoRMY8eacygUiPUjniXn2PhwEeBCp+TY5zIvx
h/mc1ofdSMIjbvxbRtqJe5gWWPkzrDY+mtSX7d9WfSmdtSFNCbIrcLDR+ZQK8ZsEJFe5GO5Edr5w
AiR/zv/v71U99qIvhlUWprAfRxO1r+GP1wNtXSWIfbzX9NCBa/pomCrwO4O5VfWObyuzaB9KiHU2
WVTuS/uky4rDyMygdWr4d510ZvQtT0EyJFukpsG2yfkOUjoYDgLTZ9xUo68GwNW4R/bK8dvD/ekb
IzIH/68za5e4wGfSl0aeruIdLwS4brqFvc3fYQiPWb0tp8my+lCm3ybhY8hzwYPQjFBaoTySqVC9
hbkyRXHBEAYLn4Eocu03EQXWJcRIOR016hPFEgmrk2eMh/TC+S3gFx5UR12Nt5qAQ3ZHiz9K6dhI
cYfAIyx4A1BuJc1Psk5GflZbRFKXr7cBgD0jRMxgE4oi6oD4WRnrsJn1Oq2GneqUEhGTBgMiZYSS
Tr38isbPqOERmNLA9tIftkf3pPE/ITaSWV6wdcMYauuaR1Qt49OoBiY4T7EUuBHY9h16/nFDw18T
WFMIJDQEVscUmeDdxZWpYUUNHhyReAUx8q56IfTeoJSsesf8E6zfcXAk/bFqcteUuFpQPc33bYdh
sAXZEifzhH/gXmBHkbmDqo7YsEyN1Wdl8kSMCSZUBHszB5Ve9eWq8DM1ugumaxLJV9lt4Zc1kKy2
ehFg1RbdyFHxykPKNwLczu66BFQcBNnjOffLxh4LwFcW6E4hgR28GsltnrMpH8AvrWkKxyGr9KEl
Pr6Bz2poDqoxLb+W3TlwmZ5riG+WCBH30hiT4HHPEcAMQIIyMoSHBtH3EX3t1hBYIJoFVUh/fKRy
ZMihOudS7SSBtiwQMn9NuUrDmdZjoxeefy27e4xm0sFhHf6fRYjzgD+kXV9FspkkQ+BJ1TNFWdge
pIVefunIn3FT6kzDWaR9KnwI5fKyhQJvDWiKia68br46cNMQW5+dPsbl02fGBz7ju+DCj4u0JiVR
oJA6nNGr+kqQEUpsJLWv8sxZNGwCUD4LB5ZmqFY3sghqOtiYsYSNgpkWgWb8weH7bc67QuCVXf2a
BLkgDNw67IB51vpP1lQshSYGGaGdqko+YvX4ajmYeabcBo8UsWg80QCcwOJZiDwHlH/EhDtkI9jD
gR3UrMiny/YZIdxHkmuGJDWCgm6ymJJl1O8zqX3ykTXlSPObzqcqfTzXl4fZglG1oRoqLfCnJFI4
wBrs9eJLnB3ciPKjns1YokppDc8Eema4OUlyLDKH1yZYGEPaXvorQg0sR0KcrVmwf9Kg68Ml30xz
2b8dUbxLn0CqXwMloNkdhs95Uz75hJKdZsZmd9m89fbf1ktcWlhHHpLNGCYQxKWK0JdOB90rNdlZ
bKSEgkAqG+qK8X1Y9d/t9R/wd3eJxEd6yMIxk/0KBBFb5zGg6J/7IcydSiU2yX6WlDJz3XGWES+P
Yp6UFkBTfDIdzxAiitbMzQYJoS5p4PtIYu2wTjjWURdGCL02sxMCkBxYJA7KuZUCz1my8pSE/ewe
YwtHstqTCjP3HIyHPaBjPsCT3ZIjVmvc8V8fW6j98zAhOloceJrq894j4VvHnsDRKAEq1tXlugB8
6b8AxJ33jYT5qXQEISQGSw8hdvpMY2AYMjagoKeVvA8O4mePtHCEm6GEac4oP7M2pm8LzO7nUilB
jnrzxdzjuHfDMhqcu0//R9/E65AC7MSL/6VEbfqnhGaZX0YKw5GA8dS/0NxwnaOusDlVgfLTiSvX
IWpGK7jhoiQ0CJWSQbLFTCOv2yyjJcwcuZkkH0F9adLjyGvRa+/OL1GcEyH4rRDtUH/QXjhQGMrb
LsyYWJuo76eCpDT40LzcsqkXewH8WXipPj/2E1FE3sGbZThay2+mzEPEomVWNxlqM4MeXclR/eDp
vrxHVTEe3NMspzZ7MIohHY9f1QoM/v2GRoFFVMq+oLgWDeGuTFhx2SUSJm3zodPBRiR5sthywOGC
DT6gyEQzo1VcqkjUaff38SGoU6QlAYYya540SGqZmqtZjDAir+W7j5bd1StL99NqmQ4uCUH1Qqee
jd92Aoka1YLX9o9xuOC74xaoKY1ufH1xVCHAgi0gYicMN0ukCfqdm8v2PhdyPi0qZRaJmPR5gR4c
QV74k/dTEQ828IcK7+fS5+ro9OXtZBk68kUdDQTBw6m8Kt9J2CEZ2S0C5h088Qqdk97PrrtxLTxl
4fNhxa01ZN8kl7qZ/OePtplDiHf+NZBJK1EWBLNWbgeexVrHYS/JUraE27GCkAmlWsSbMXr0NXL6
Jkkb/AkiTheR4HgKfl/OKmcVyqTYmJAHTikPd6af+vY0d7kp2tJvCZkvr5vgPdndCxWD+NcA7KlX
RpU+q4CvVLMp4WaKNkMpBCNkv6JTNsuGhcLNQlG9z6OdzAcMdtiRbeGHJ0Hw9tWsVse05FcZUcZO
8IhvWm9OW/zEYeccDhoWXwYdMuPUgxhhaeN9au+Q2RLcQBt9BaXcQ13u4iBxmO3qTmpx5FinWY0s
IPR8AaBUjWbnsrLsMIgIUxTDb0bXuHvumkh9xwDgeXa9Lzcd5R18TGoQelhj4OZ7d6OG5txTnR5l
WzKRSSUNGRlPc/wkduawfUlPCScEhT9+puZiq+QerrJjvMDW1zi5dlg9ymrf7vxS4FN6bYHZpuvW
rXn7bpPPgPR7fztsM+6RqwHzcllGLnrryuvSZ/0iEUMxNlAEPMHkhrjUDy74HF/YsgPvdedyP4Xg
Nfjy1Ja2vJmd5B2SYhZvhMKqPhxu1kaZLR3kEis6j4dqfXqyNNnJzJMf2AFYknaRCUutmbFl8DTI
8mYGejt9XMmlqAK268BVgIO3R/WW22BisoznRDSacKTDk0/q0ybxKL2i7OJ0l3dxZhmjS0pVAz6D
8kq6ogq8zWg83FRy51odr25294g7CTLGqazfqIzxJpx3et7i4GnCe017zf3d9np8mFYzYgIOB89X
qPmEWfbGGbCBL2o5OCtkWz80BKBCOHeCKXRW99EJU9Avevk0l8r2O4z4ie71YI3FqtOYLl0I/7L8
mo6CEd7Nv1FK7C0OgeDK7mYuW2pnZjC7CuP8Gdr3h3alL6SesQWbppQGC9f6cHG+Gh0R0WjyOYKc
OCn0DFu0KbvKUtCGTBYa10C6nPpVy/Jr8QuSsAcNodkHCKpccoRzbD0HDeMLfK1zQgg7jY/YIu5q
1HBKcB9C1sctdcB6rqi9AbLmvisFaiMCGXxgQ62GKG9SEx4qoh3xVqoYmJBIVvb29LikytQiKsyj
i6bf064NqFTqZy0Q9RglvzugtBZLIVGuqDEn9QJbYFpzUxuz3SBmkgX71PNqAmZgRLZxySM1+vhw
DXLobE4ugzQVMEqDNbMcKS+KtUQK4BW55tYxl3oQOpcQkoh8VJHyNtU7KzWTTdoW9VZ9ms5jc5ii
l1kGYmvFNDFLLHxfsFiTgCHd+IJiXAhMK5AtJAn6XNcMPGdRItJUyErjUPSi1OuG0gUmn0kgWhJa
qS/vNZVqIOAyCxYUskH54DKtJPlBqZo5vHQlcxf+JMJaNY+tbsEVYyj0F3UKCIOTBMC7y+DtGpva
lFqV/6W1zQiFsuT1EHiu35Nlcztg6kn5PnB1imnF5rNpF8gMhHEsHGGn8YiABfS3vzta7otEXcmR
CJPG8RqeI9La2TAMwlZ+VgJiVHDGqJJPzR9WiCrW0uTOC2k34AFhTHyhBzi6AkCYAM5xtH4B32/n
VqXL+cu0SCqNhksaSlF9bq+OWML9/P5dWIuXB6eB89hd40RkpUlrd+bGRG/yNiuERBQK63h8UkYE
XORUFd/Keleogs6ccPXKBejVlU+G/acPdVTziPn5DvW6AyRS7YnqiDUX31/20SLJBNCop4Y/+BLG
b/UfTk0Xh/g3ah/ZDy7cjjjJmVICoYUZFfX/ZLwlHJMH3eLaNY1thzv8cypWsIUsB2YGq0qhooVk
Jq0McACbiqyjAcCQ/UVWMCz2O29vjqgFpxFw2QHgtDpq2n8SbTvEhJTvtG/wcK23eGsgAnwL30DH
yE5KglxPlkBgZlF8jrZIALqowdmw4K+xpg0y1Ib6b9HMtTS+vFEJ1J0IFsGOr5BgXR3gVcCgBgLc
iDFICKAkvCYHvqjfOP94mQB5b2RRrYslSHwO5jHdXNCqdIFyoU9nt9/l6bZoB7SjK2+fhM3DkjHg
ANBTZzBdA9mI3QbVkJDC0jZWJB5wbIYuFyStQLrkZrxAOooyO1nrlpvM4RMEgok2TA2BWRhx8DHF
rUW7Rz+r1BzAcsYqgOyfPZXtakw3MstqEpxeVmis29RAp0YFqpzTIN40h9GALW9lopp+z8s43aas
SonEhZA9osT0mSw24kLd3nxVlnOE9JaMsUcrpX3frFpxU29GqqcOi/Y4JQV5USVYQKPrKdVqdQ96
SnS71S7oV1gep4+KsVWODKj9M3lXHQQNCeCuwL3EMofWzFR5NmdRSGw3fJXASM8kyWFwQF+VQdef
JxbzzBtUhZpK92r1jQKgbcZbWLYAGGVNgEg5KJdUz/y1cgU//1NdcuftETMSjFyPQmW1taODwbWV
/hNp9hDCjrHAWv/KtMwEHTS1tLNzpcw6tppoE7aAbWag7Dt0AF+6XGx8JRokrfpfswuR00DXv0d1
vOP/U2v6z0ppZwAPe51U/gRdHCCweUC98iaW8NPml6WG9It94D7qypn+6KKkultmamlUVYkMlCYo
cBrZT82auoVMjNx9HXZAxDPV9tvcA/p6vcRGuC4dwKlXhbSG2Wa2KkKDUSjQFvNVHjSjBWh/5Tui
XcpueQn7hnTnkuUnK1H6NaAfmy4mz+kjWQZT3Jr7cUdTs4EFupGVUzyHM5/ZkVMPs3YVQrLI4a4Q
61ZcTMUY95Aad2XYoBGC0yRJGToGcOAnvspWfHDtjvImN1pqpEKOouspfTEBHVRQW5G1WP4h6ehN
Ol2eMLwd/GsOY++FSlcxavzOtODP7+MoELe++YUs5OZNTYhdpg8y/jvvYXdnzXhLZ6bfRmzJzuKx
1SWuPt6zxxdpf2F4cf/iWZKzoNH1BCL6bFS8tsca+0WbGqIxtZ679/PpqHOsDYIhNl2YpIP8L53h
nJ1scPO/iggrKRl9Zvmg09U7TPNO74tSXw9oPrX5qYlapDxypBGu41gX0IEH1b6KEbWZcyHvSLS3
036gwGCTExwPpc3io5FP4pu1Scu+B4Sw8Me/baCt5hgBK0t5yaWMbQIHhd/ncgRTGdk+1SBbolVc
6vlbxtvDdgQPZb+FzkPl9q4dfmQk01RCkELS6PYzjmKpqdPWfkYi8qFHfF39KUJV8BYIAn2zqYz1
Cg+8hrqHwwgXbKBGiyXc3VhAX2T0tsKYlPFPLQfmEOkXd4BuC5jyDLfmR/YUV/CcBxwI6PgIJsER
3YUv/GB0S5adrwdI84453e2MUiGusmdw5pDQirRL74bT1ECPsIEyN7MC5CphMACvFnnXr0OY9wHZ
QR7eongu0gG6BWLCTx7Kffg5sOs6Tcux79NVTtD7tyUg+VyCcO/z0l5cuZMD/2hAyVKbJ0VFo9Mq
kwuads45/MpKWr+s7WX1xrNQyAJR/TTtYoRG7dalX7UQYV5u9l57ZTYsgAXIzZKyuQsJ1tq+TNx5
DLuPpwyBjuwEKQ7bdGPHMK80hyh4GXILF9GXfCpxCTDFUa2Vz7Quw1CbnCAnDAJHda4EpHImxdKB
QBDi2QnDpaSmqHKUqQaMFklq2z93QaRQ018i3gyAcxiG45gkO4xwsyg49NAlDJoMNrXk8w6CiRSU
PDo6Aw41iUmSBl2+xSYLouCSz4pXcksIIr9JUFRPncOEg0sTj9hqsWVtQ4dLtaaNuM7fSAo/qv1o
PelM6EpJ8w7rtQahejLQ8iEr3OrM3kUJoTqTFJkJWfUFUXa6DP0ZX5Xkoan1cUcgN5kSg+yAYT68
TtSrz9plPy1CHpagJe9Uv7FnMqY+QGbGAPQaVHDhDZ1sFD5Vp5JsURbiDth7+e8pMqTHXVYCPzdV
avInwCB1YOllsS3bxCygKrln6bPjKC/hMlqjRBltCj+i/o0CcHNJ69bNpL4CaU2O+AGA2ZRsPhI5
LK4SIkweUr1C3I8MJTGuEsK9pcUBgKDkVfp1MS7ouLEoN+oSy9yjeuUb2i/ne8kdrTWnaIeQHZV3
CIOALWpRTyWqRuMC7PbOjD3UIm7VcHI04X6+KhHsorZAeQeli+VCRZ0Cvi2vEjbYsKAF4NL5EWjg
UODi7gjmAtdGBsZFLKbLGPi11xdjLsF4VHBpiYMEcwHGPMT7hP2EqaOQwDZFzJ5eg5uYzZ3AnYa7
vPeDaYdUEfOZq1J3/7ssBRPGKwW4zu//4BZGPPtggZNxwBMIpY4GSikHmJrGDuCZ2vTo20vcfF/0
Ms0qBiu8QpH43G3Q71kUM5O1DGvWdGPfaWZkv2+oxHl4Rjm2EU5ZBUOLmAwgjJN7PHAKlt/i/OL3
WFs+kG53rR/MQhLcpuKD0xkh3jItiEfqqWer6PJ3BZGKMuQdMazDQezb8f/D7qg0eBaDk9Ucp6z2
yCthE707Aum15bvunmHVqsmwap5vhYFeUctl4YeA65tL18D5TKrW+RxtXyRjrSWMy1YzbLA4qLrU
Xg9ELizsx8JBWEurohRWPg7xelRpfHd+LFrmmU+iKvRF6jPyl1Ud5zTMd3ixQ8+DRytcgibWocL0
ASyi2dhVMk1JohToAhEiEx/jQroMbcVzC+pE6un5bhOGnXVZeLJVWa6Pb/I4E2yPslbYYiOATy2v
rPhEsLPYoHpaaTtKJlhHMbMGSPsoZ9ulIL74iQZ5WlGkvWpBQhJM2LdzbqXn3e3r7+dSxQG8UbyT
vuhFUguOG3OpW86Kdu2RAe0KtmNTYtnYgSBgDTzjK+Rqkrkg0bhP8OuDXSlTuFoqMwHOGeyv2fnv
mPHTV2XiQp3bcLE9kW4QpBaAzc9l0oZK8zw+wJRNyJXuOb+/nm77lmApMM4NFKi8YBb5lPaiv+zp
T7be2mlQbwi0TgphUhwPAMyVwzwjBx4HQQMPEu6lPYdeWIPkpOda+7Ge9g4Pj0402os3dF+g6epO
W5tz4qDJWYhnZNzSl8W2BpcDj9Thkf2saVb4hZrtsvJypm+7/YjWVHOEXBdLiY32MhpUefFlzCPS
EB17/dXg5e7ZYaAanDQcrkyvHn8dXIT7L5MOVVoyiqWpj1TSONmRFP357rvpj5uguV2V0kdapxaF
PD6WR88toOQZIJ3x1rF+efmnrLWIWBvA4IKq43mMEUhtKw5054cTyTrGM9CMeQJwUEPF6Vc5QbQk
VQr/92knzH2IBdgfZUZw/34Q+GGtJj0m+zCK/9InGys4qG+nAYFgnIjN0eRtrdgboUqKOEzlxpPN
Me0eszaTv5re1Dv6TGNNIJPRRygBcS2dcBVeyc+3RULjpiVMXx50jX7DF5BNJfb9Wn6KTFCVbP3+
dib/8mPBDI8hr2dzQRpUUhKPGSCx+BArdk4lKqERxLCRz6sX7mMPc12GxejpHo/ftBjzcT1TMFqb
Nd2OnZVeq5kXRwfgcfnjn9zwYuSj8r/wwrWmQTiV7PU7nvXmeAZkKnUrIu+gvZqP3W3Mz2q6bygm
ylFD2Z6dWyUvUJtfaQII/QiHzo1TZXUhuPQFQ/U95j5ePuMFa6gqE8sbiaODy2I5fC99bV+NEnBS
GOOX167vspAbetLTBE3skmhOAA9zTjtXEboYKffHKAxzb3vtVJHgWyeR1ISHRq35sSZszsNKNyFF
rBkGVuE/k7kqkynDGrwO8KLjgTFNRL6yYnJLOI0slW9DLmMZMq3GPnU6DDbKBMTIV9jHnkZU44Dw
rUHAdRhvw7bCknvZkaVcpEfsRiLucj47apmN2GvGiC6s4fj0xKBRnbE0LDuyAZgI404ZtRUSIE+q
BwFTRRIuilCxkvtLghxAdMzQRqXQ/Q9sNSbq1dvbpxR8jVjkfLLQtWmU9QYtFTupezipZSW3Tn3s
Bspn+6CkJS9BZpzYlSRDTp8ghggc4EnZN//ZRc+S+aSfuQUN3+JogtlMtDA3zcm8NPmBhuBDKUKl
jYRmIr3igEpMiXM4jnOg3T3rbqexaNZzbRAwxPoQ9sTbjxIwWYpHEaa0YyzUWGZ5rG3nBwQs0NUQ
S80tgbGT0VJOb5mc4QmIg3QtP4gm4+xIgBkpvRKzbPxsixRpoI1QCthxFtudYl4MCyh4ETU0ZBhf
boiSUW4shN7BzsOW8ckaTH+R9tieAUM5lOb6SXqnjGwbAyMSzskwZxWJDb5p3M1XxQq7aDUhbAUD
meeD2QToaVQymedKCtPHtvnSKBEpHZrJn4eTUVWU60BHPnpYEGooCBYeH65dStodCkBujlztAhaN
vSob3QZOomitv2TVRJ9QJlUkbPiujic2lwV6aomXxIJ4ZVeVmzSn33Qza3BpDH8fSbYx+bIuU2he
gFMa7OV8bEQYVjYH8WxpBdDhGcYJ32+3yehgVYyGTng1Euqfph5OepIFGkfvYOtgiQzJtIKOc1IJ
MaWQcalLb80Xe5fXH48buc8noAUZ1hyqk9AtvEYtBxmE4TUyHK1ovUtIrSHzmq0G9CmPU+geyCjp
urxGXe+38l4izuRi1akTypvzhJw/ed7/MjayNAdnyb9MwsR0Z0RyO2FTggNe6wo0ZqqviG982Y6f
5zlhuH5Y4bwc0Q8kLW16/Lmhm04vYypzw0XNjLHES5wNWy48UEh4EGExK7Y4ZMnzxco0zPidblWC
tRtG8v/669RGBVB1VstpI4KNnll9KkE0ArjZ5//WNZxj4z5/MHdH5oEq6hsJakNRpqr9fK+mC7GZ
XPnNQGRBIv0Rp6RSrXlyBIugfPOwE7w+gbQqhr8vLiPfaOqo5MS3qkbmVrNkjgQXBRwOU97A+zwn
GUIH9jlgA9GJh3x3L1JzfJm04L2zFpvXBLo7WkMB6HqPGglSX4IkiUJolNBRncJjrZpIB/4BRffs
hxfrgWrz2VN50tkQoifBFH4SxTYFQPrsyfO4kzqeIcmSj9W6VjXxFzHNqS/q0IqL39l3t12Beh49
HwIcAcWC80V499R1q+o1i3b08fkXf8wjTmururaAHNCbPUfdEamWADrkTR/IAiqlhJYb2Ng9AbeI
M9zUobe74IKFKH41KFlK31Jg1aF8PGgZySxG1CFRQ3MxvhPKA02C5VRZMQWxyMBnnb4xSMOdWryH
9Pg0rc77yon7vjP+i3FnFoopsEqQPS2v0hhZi7e2HaKnFg2NNYhl1AcAdkRTgcpE21P3HsvOmnjQ
w2s6r9i30j5wQallMwEibAenhb58SoiA7oG/dii+DzLOEaC2AiWldKL+V1avkNthkUYJ66QbqEsj
Q0ll8PKTXkodC2Pu19lFUjH4sXKqr+YpHuhij3P0l7VSl6ZHMMgqLisxolyIVofP6v7D8XGG5BD5
yePjfKjRUjrJClb6Q53Lr1k4pF6ZqIvt9gvW+dGeFJIstOhWw0d3h72rNOo/xWki9iAlBgM74kE7
g1yw9Wx/ILcEjbVp/KsQWKyCTDa3WoGDKHylYWQ813DVaUxSipuKBrUrLHcZNjYjDUqtLSugDrjx
N5spnstWSYM6VNO5W5MR8qZJ+85vDhCFFHK0+MJanyXIPpwhY1K5DlLs5WTYf2ZKxBBxwayPAFee
t1C+f5R9axD+DypFG+2dvZF0U1EX257F/RvZ4GYYvauYPDwIMhY9sJkyVhZeW3RR5GUxvvPEKaKq
9Coa5BTNWHRjSKwtb15CK6JG4mry5a5hszIU4OkN485Ni32Cbo4QVlzvfNyO2syefuUdbKUqn9/6
Z1KCNjMpJQvQslsi7J8Ks83Oy9YsBeK63LbubDNltn+KjSDnZhSbRg24x2uLZ8bVVwnN72vqo1t/
Up7Pr23UVpTVDOojaTdFu9EZVrmhzIFCXl0Ls/r8IeYJrl2k5UDCibpc2VT5qcw9goWQhMpq7xt7
Oy31j+YG9b4NyeCoHcH8vBIuR2oPh9I9oJrhGBeo2v0h7Z8pjWgy9j2lubKTp9Ri8dXJ34Y4gVOo
O9fk8XwmaGOiwhNif0IsOqORHN9xp5pe0OL1UCrW77j+xFwAkT6v8bPHLywdUpSopQPZ0/TU8s9u
KU55f54uo7f7CIlwpFO5TNA/28i1ihIZgRYJwzH6fEDs12XU8nh8oSv6uShBetBoh691+iZHnXr4
d51aCckQ93YWfh+/RaKRt0hCW669nd8dmOWa3eTdq6J0u9gkpEQjxlhKaClLRKmAfXk6JL6hVkk+
nD+2dpMzisGt/WgnynVKG/rl8q0k7aahVMjENBRNxbQRaRnqZZfJzafDU//DHWYJ8E9v40SeLyRI
btUpPBhEnGrOCml9EUOqOei7fxB7a8PxSEpkEZvlnlLvJISHIEzsGovk3FCipDbVTt3mC6T27/zM
k1OH+kqPopJ/orq1b4+5Rn+hNn8/z+rQU4/duV9d9BLu9C7cjZD/6AJwTylUmvj5eyW7K5DJr9g2
jzSlBgiYuQKW1sKEyl8C64sOZvxKWBPLQlneVmrN71605TdXQGJRMGBUI5lWmRFSX9q4kfCPMTax
RDC7KEB9vkSVfTRrjhl72MWlO8haV2hs0z76caK1uUM8Q9FJ2lFkSMfjacZA1gc+GNnRGokSzcOH
9o7En2A+lN0PrgaeqZg/d+w5R5mpVXF/Jfo15DG4nGtXR2ORhkJuPFjKhCwjekiIpk1XofFtvOim
WeVk54N1/6Gt6IwO5oZ1kXxbmKVT+tHcULufZL2P4kcM1U+2VfnZcEk/UnClLUN+B06z5v2wTiDa
BIPHgMbAvZA6Kazgh9otI6BPvXDQz3kmEq7JKU4tL3TRSCZteMTjQ5wSik4N5YVG2s0Sa2hSJj7E
4HWgMPGOXVq8jMULXrNOKvswnBh3Ovp5BnofdJqTPBnOgHQHFKLFkhILwxNbo4+fCnWXSDuRqyUV
3OsowiBmFNMEn8/12BIX2qRrZsN1jwDVX6CiTyCU+CX4xIzY6QyTTXmHSNIhTa9fJqA7ZnwCF/W9
UKSoLmmGF75ubLTzHDeOWtEJYN2cQfEzHardDh7ERmCnCC+Q9u3wDvBgCwkvdVor2Auty9BCs/9p
KYNElS9MC/KCEtJaT9y6yBCToMZL0bucdkBUFVmrmJNpIxU5UBU49Yg9Xd7YiwYrLqpD6cQklm6l
ZHKtFwVfJGhWDDRBSJbnjRxhsPTYtRf3SapCxk5tgvLs19LrhBhMFqMu5XKDBog/e2DQOnjR6ctC
Zasc5bEOBFwXhfgpkE4eD6DwSSUZ4TMvzRatyVhK1VQa7vo4BgpfoH+nm9cr0iZtcuIhBYzCksyO
70ZjG6ypAulwBr6AF1FhC9ZJJPh0sh1ysIen3S+pGDGd7fXqa8YzhYOa2vYgVXCYgkao6jroUUjs
XPhB2pABHszbH6IwsK2W48c54S9GxIoW/l/un2Dpp1Lr9D5teyqzy6OlU5eX2FoAL4xKmBO1j1qD
tDtM2UkZpaPfSdiu2hnJBXuZ1qf3x6TJeWZtYeHtn7AwJ6bsxkROV76WeQxV0SAr6mO4uRhucTWQ
aX80UHj3qewBQr3uOxVIYkbsTuOG1JRs7BZYPsrUTRCSvBia+S9A5QRvmQsJUWQbMSDgiFhY2M7x
EF5X7mZooC29JWWaghURih8aCmou6X9hGe+bct3k6qiN4laQYsiBYiourX2XkGjIG7inlUxxTOXq
al9OWMDhZbFvS8SA6JLJO3M31hlwT4OCVAWngeWv3dV+YyU95OYt3pYFt2x75nn8N3KmxlfHp24b
CZvbwApOvOQPDWTCTh3M7av/tuV50/r/7Y9Uw4FNdVfzfqNi+rIC6HYQXugwU3surZcVI3yuCVV8
T+y/O49nXtyhz6Pi4JsQEFg1PDcw6dVTkLTMjVKUz6eleG+xyhKfuL8AkfoTSeXZxNQrPjEEMijq
pz5y4QqXL7qfdIJgZui1IAOpp03mXwgRKlvpub4Ho7k8p5fbeKrI41wCyQWy8cIxP9Zs48BaXt9R
R0toP4yEEvXrip+FQdYHsBUxmOwqeMz1Iv7GUs1louwnRW3MyBNo9OZmc1Gn+VBVg4srvyRc1OZs
C75WForfgXt71t9jLEdGDQribl48hTc3TF7VPycRTcOoQeEljq5jXz+tUC2pjm3q0R6l7VjYajJ9
ulL2xYxhs2yvBqpLsBwUmOqrzxZATnt6eIi4rmQAr8mZ2o7fVbJl7dS1ODucq//6YXioZRQ5YRSd
ruQrcuUZQpPbkn/6mkTZomnu4v8G5vW8YkZ5NlBb3UkuEy/hc4X5Bf6JQ++wMj3GbBe5IgawR93Q
E0GBlx43UNNpLPHZDeRWW8YIlvZjKodZ+OXjv8RaHGQrJLLBMGdTqIrEHcgTdGJKLz8hCRQdKJg7
j5AFWHb+9KQtoEPJr3DrIT7jNDubU5F5Gxz06dEGVwTbiyihTuQDAqoiWF/qlm9ibkTI65KBxQCM
0BL/j8393iD62RHMwBxXlQZtycuxwdZzTbjEReLDIIbNn0qgQqc14qYN/MamgYiH1DN+o2c593UG
CirP1cL2V47QaIiFiGuMeNG55cwSX4lGoiFEiastcF0yP8CIPn4MjrBQAjQMnFC+7w3O8hAgLnrA
/F/xJIrwA2OFhtMjOARMibgiU04+0Am6coU2xEJjidBV66jvAvSYgXWw+0dO+bZK/bsafHt7Yeto
noFOJiTacNy/LcAyj+8YtJAnn4HO8qfomuHRAfThZIJUxl+WHKl6c6dlXZWed4tkMOHhmQGSy3dh
eM9Rt4jNWr6zIoiTygovRm79yCxgcOWpMug01uhTf/wxOn+3Khq2tWdU2y/TfTXlgmxI66OCBcV/
qjGWmAkhxs7Q3np/rh8Dp1YloMP99fWDjgOaxvvgWlz1hxigyHiolBsoVrUM6QDCAjAyHhBLrzha
QJlqlVNqnB3rxNHYQuTF6EJL6lAgVZLwMRvtL+2GTssN9NXaJLX3cTuLy7XjrGT3tTW7TWVGU4yf
EI5CZseM21VSUxAYXZUhTZkDAH6B7SL2qkjZitZdlU0/q+rJtCoN+jRKj/kEvvSop+07IGQZPZQq
ik75TLBxD1fvI26vY6EVLrnQnf5WvUdBnZkd5sPJFZWwCsyD3rnuNOd6v9qaQya4D9tlp3s54jPx
2l8WFUPtrpBWhcR8mL13LtQqP1mhKNyc0ONQTOITNqF8Gr6nW6O0QzY+Vz4pSXqYSSfGP0pcYb1k
Smluid4DfsPIJ7vP87qVgAtauCbSLQfx0cYdWniRBKUyJAX4wz78xzjgO2n67HBearAx6b0HefUJ
R6A6s4LZ/Hz3i6ny+HujevBeSUDQEx8vA0jutLLhkVvx8XXdKmYlvi/vT/k1+Xk3J3pN67BfHSxl
nz8gZj3GMpltsZ9XVcRrAEI0DMPutPaKRU/STH/QFNWBZa4SY4wyIR52UWHDpUgM5aMC+b91H0Z4
8LW4tfr8xjEIk2NOaWQZVI2j8dru3Qak1WpjcbJ7kGT0LYJZJHwmwsPEenSBSPCa3MSL3FZCYE+b
2TKFZfb2bowJOKSOQ2lsbz9xsS6+VnvDsSynrLi/C16mfEiAUNxrh/8RgZJl+NN9Q9TpvV2qdUr+
M3mrgbABjdAUUyt5Ir07yLpwlAri4o0wniMc4sezjPHosMPy8UouejTlHfoXHUiAqq0LO0e//mQv
Oszh4am2lvcmgXwY/iYzizZ6Si/KDsvVQC0Sh9fc9EY/dT2+akx8knFS3SuLptCTfMKCYxmkMW4s
cLYS17Zo2HTC2zzmRL+VCm75zVpwtvOCR+4hKHATTPAKf5NrIN/ejAj84r34SwxxGHRnREUBwerM
oxhu7rUTqd4OJPE69m8vM0UiJKaUxCVSWpCUNzWTXQofgsIzE+TbKSr/BL/JCV6rFbBZWowDiM4C
VkKjtMtN0wpfQBeifkiioIOBsvw1iE6cWpWHBywc2f79QYu6VERQAOxiX2a6opxCC+5kFz4kCT0P
A2aEjXO6R2rFwjqoKa4ucTlGzTxVXIK+GZX0j9t3vZ5++rPUArA3wht/okF/rs0y+H8Kf+8AXx5u
LGSVKJzkzeaJhYyHAWQw5+DNmKPIWRBcFqXRdVet+AeW2OKyz5x3mxmzuWKWHZXpVjeQsgb+aTnD
pp6sy8Gf3hKkcsOa8+gGLkGxL+aE22/4DmRVFnquDB3993ABu2AWeow+UKFwdMF7wKb57Odc8nVY
76e1yCTNhY0LXMVXM5zZpIHngJXsPzJYKKlMYw+Oc4GZz1PbJ4OX+ZUz+5PoUTefUQKQiP6ME8uQ
/JRsOKNFldOZCvGtjuw05WeTcGSsiZlVHX4Tx6uXEIUQWkCeI6BixAL2lSaT29BiDlAo6RvDoxeP
htQO2McFWKle2CIf0SmWtbTgRuSPvm+BDi/PN4RtArvsl/FDl3LGYKt9Og0AAMDOVx71k5XH//Dg
Gskv4HFU9XrJE2PKxAdvrVBC1VhP8SubuaxyL5rIrsvaipexKUX7QHJoXK13GW9BV+nAs2OSeGp3
tEp7cJCL62mQXjIK/G6FJkaNQ9UG/lpXvgrkFKASh7tD9IHqc/XU2l1fQuY23H9CBSlrJZ2WnGil
8CLYn2obSe/uUnfmxR3cumgwuB4QFo6cbNhutesla+RZ5mfPpzUyxQlaDOFotxXrMwAywjap9f2A
JsREG+fnVtB6leGfMZifkCaiQX9VnMZwGW4Gx5OQZ1rXxluPSJd+E4r3IuZAAvd6Rfk7NFMyOXQ9
xn9pd2fzuJCxOfQitTPNvl8b8b5XQgvBlfSJugCon3X4npgrz9hAoDZQa2F1M/3Emb2lZBQ0rwE/
JKS3FKee5st1pE9TtS3dVPw4JCgmQEsB0ukRTnY1RDGXtOzgqGqtYiAzComouuUngWCL+6KFJTNr
fUmNGHKcS7SBAnFHGkzXIHkCTW01wOV+oeE6272bDk9K/3LT54iNfWwawxITs08nus6ozF/2RvZQ
qS+Op4EJcT0iuA04OmDp+Hqkwp8bLFNzBsk1S22+Fs4CZkNHA0VgTAjkLfuDTSwn+4t3+cEvDMRD
IQIH5qQMheFJguwuXTK/UHKFrgNEM+pY/Yv/aeCSL9BTAzaVFyEaTSxMJO9oEm5u20m87YeMR4OY
68RCgn/AhQFPsP2J30Jp6zfhxGzHb7tcw6cd6dt3oARis+MufpndZynrY34u3Kroro4pcymOGHHl
3Rf3JnVcoj7tDIIBfNxKSPfTcuKs4y65Io7+pdX5tU7oyQHAmc5LtVrmAp3B/A5tZ0EtRrmQimWo
A+9O//aQlXOw29l1BJKVJb0hlUes8mtAhHH6iKjFhB0KH8gezGZqykp8GKpxDXd/Muql39wlNUUT
PShoL2jpbDjyRaPNExNQMDl8g8G8iGtHQ6GYVLLJbLoGyZxBasAlUpc2nVYtnC6RybS4lzAKFiy1
f3tkkyoPfG6QBR3XElia766Ab+FEEbhNuhufvhVUPig6sctW4iK1MPbGeSJ/fc19wbz2DUVvzlST
iZ/SsOmEpkbDA1N166FU/l7+mseAwqoYDEeT9l5O7XxWIOILEH8cKO433nk8W0NN046gdJff1k/L
MZNhcowepCcHYc3P7d7LPXvODssePu28Vw+Z5CIGxfWk8NOtQzKtYiHnZJ0p9G7DFgVHYAgCtCeQ
ilMAPqwTD+BEBYyep8hZNEDWLcy6jiYPtNohO6dVVBr9ER0LEmQygODCog3ogxJlaqG86hiYZZHo
4w14UFC5KQ/6j0XMPXauedKDkIYqsD9D67gCrYekJ4C8BmyioHlXPWIxKnLiSU83Yx8y2LRuHwDB
FPk3IZvE3YXxCZWOppdra3U8QocoLDglLletiIvGmzhM3GY/NuNxpvk8eOhVaPqlugrms83at2Wp
TRgS1PDrjhnL3KT6Muk038O692vtuvEB1AG0R2SLsNY7A2Y6pI8DCftlb0EgTZkn/sVRX5DYig/C
2eVjzJ805m/YdApAA5F06hqnmLyQfuQe2vHNpaOni+tIWttI3DGoChIUMiFxNxRvW3ocVczh0tUp
amwu3rkM3gO2UfWChAktQhrmfc2Nh/c2g1gs+bZM8rPUUE3rAkOXjlkdEBlejmlIRKAni5DgUbt6
f0T2KuC2wg+MzFq8fQzAuPL0lhKgErNTd+ucEelECQVSaWNkctOoXRqRIXkcECJ4WU6EycPrj5BQ
LUYAsVImWkvQyRl8DFAwznRcOYHf+84P8So+cAVvH2TaeQezQyUTTjtDGVt6lLstLq7ogKyujUUJ
Yb5VgSg28QJtzlhodmY1ATDBqVFa9Q+fjEk7mI6c6jUQzH/W1AQg3vAi9Xkd2jhdafvAUUC+uu+8
v59yfNSk51ZgMXR+9ufeN5Yh0wfZ8Agze54Syst8qpwgC8WuFN+uclTktaD9EUClhAcqyx6ZYu4t
Rlwe7aCpM3uvZ4Sd4xUrpXLYUkOUvrHwXFtBwVNcrsC991rGbxoWAKn64QmlWfo1RJgcFSHNl7K4
MZhTVAz2SN0yTm8UQocUkPHgKo1G2ONQAt5ZL3uDgZ8iiIcHj1xRSWzeVAWDGEjreNIcp+1GcUHu
DQRG2gLO2+U7mBbQ39d2jclnaAPkJAHbNddBgqTw93JKzhO5QFKwRMiDIZOVPmEYXKRz1EBCvFJQ
9AxjlECViPzGHhxWygb0qP/lOSPIob/9wSq0yCJaEXhMitGwQ791iNv63Hl47bmO1UWN3yIPcHSr
RurpfRKmIWjpmYFaE9+XJHVEgEf/0651ZoxSocaMt9Bup3xeEVJmU9wCuVM4THc6CqpYAvvt6CoA
sSNRSveVLEx5OyBYbxKAtMZEBipvB0RfyxRTeGdxvqg/tenn5S/+uq5i0LUin3Uepxqbd2oOSXxT
Huqe6CYYojjX34I9lQ1KnC2jn+gsVRP8E8kxlUCicv7gVG5+31EvH+xXculsi645uv637v/fgm3F
XH+I4x5O2ZkQmoFent9HhjvlzehU3C1r0CD9pgxSDhPotl2YYhibSD3TRoN2P3+cHcnRUaLkPQbz
fWVR3/YPJI1cn/VfGjPzNSWcB9NfREQrWH3JZr+OuXkmx62sUjDLQC9Ej3LCqew9rSitrdJuo+yf
ea4kkMDkZnlzRyjhfm3ul1ULaCgAWYpXQUZyovDsg65RgZ4rZBAy5WzMmSr9Z/u1Y0QdDP1xgpsv
UqCOi7glbJAhGhavIe+2O9ZdhrN5jOm5DNk0M15jU5LZw0e7NNbeKHBhwGj/2Whv2uIsXBW3MCOv
55DpeSophcA6+1AqrR1XjRPKrDEH6o6zh7L03enqKhKW4+ZujwjC/xZGtnFZLB6dxdnX1h4an9yX
cRZU5uXreI6nXsWkiNWIcgL8aZnn0+UhEud7fPP7nPGazqGoIb4SKdvrAOQZyF6MTgnpSQyNeNhA
hRi/JdcuFOcIwVIUp7JpzecO1cKRRRTOsseZj3vpAXXz8XPYJII6NXqoxBJtFseT5nQdM3OTrDJh
Fm47ex3gW3a7K+1AiIjyHGWKFbiBPiQeWJE8zjsJRsajfr7mop9dCKkNh0UZVTMEttQATIIG5oY8
GEWluOTiL2c1oUWjGIlkTBMGH+VMSY5QtIu5/i+WEwS8mhiLlb82F1FnVPKB+wxLJkREwsBukV7e
apIjDJRg1GPTaxV8Hsch135EV174bgcQ3uS7EHBHWTUc9r7Puix3y+MnlbBfdcCcg4n6W/ZRLK3l
MXT+T0UKCW5eNXsOnyxOF6Lzs54hxH/FzuFYlQxwKHpyPr32Vg/cEnZ1NTutf/ToDPVXPJRmSBK9
1DzA2Q7cuzTrGWOkCPcdTLx+uqE0fQkXVF8RamenBgi3eqrqTEOULgLARhtrUEFC5DqVTEqAnZzb
4xelA+qrTS/95rKuON7YJpsL7+XteXd/A51rxEFc/jTZFGL6+Z+S8Zx1cfy+d5P8SodJnFKx4Ygz
LZLpgF5r7Fl0Y85rx3BGIucyTN3OKqVi3DgT9PQP/kRDA0YUzLn2SuVoT5QavLfxWsTwW79sZIBl
3VBtK8nhcrsAICguXUy08bdZRwJSHDsiVMdebQgatozTFtXYud8w4rZKAICOJZKZHQCJwrNM59E6
5tm8R1RsU6SPZcegcr9tc3x567nVIU3JsyqZg7YhiF8LAYIkIi/YKwaUPgBqn7CTlIoHhTyW1J40
vPkTgaMcfrkmihSMkvi0XGpJHcCRhIDT4wAWpuwSLc59rQKgN6JJLtDe089izMe61j/xQlyUPaJQ
6K6VKdZITauNYITmkGgY3droev3YjqEjmhvGptgV/wIKJD2CZiORy/d+B3z1VOGs679Tz6x/NFh6
opGMIqMvPaN6Mbxkg18TGicZ4GkbcUdjWEcs5SnXYmmz2ruKAa5C+oDgU/crD1B+9oqGjpkPtmdz
csHcOYSXScAToaVc4fgkPZ0rSTgCiCOzVr3muACeg/4OqrFmGvVDIYJ6z9WnFzRIW/3TQWBQGdan
EllGUhefxVphi72ZiiPx8TuM+I5KxxSNYc6gy//DJqPfwwuW6SdJbLlxAhbt1vQIrBiLLjv33gl9
Cqsx3ZN9QADIXnZB5pXfIqncuwvzso5gg4YeRP0jcrZVGCVqLpCT/y4sPW3SSMYXsdx83Xd1WhPs
FxuGS4wAnJT0mdvqXGOFRgJfWGYWbqp4+D2W101P+89zSveVZ/oeTkx2dNyAOq/ZZXBcHoSw30r8
k2bMVfByEYajOmCBWfVYIN2ChxJkuWHwpLjg9aR7aVu2ZzSRa/EJog1icWMVyhIYFg40ESPWmc5z
92TMV0+LlPIMA4MvUKm7zPy7fCJ4xjmiU6zIBCXApSoJwY5YAfdkVZcF0y8ZGkSr3IOGw5rd8/Xu
jNDBJpPY+Pu2Ms17GZIdCrm6gaLPC8R/sG0medvCUi+iPpHNCT+3UO/H64g2tgr8lEX59LzryWDB
V5OmgrDqYVzAZ84y1Zk7urKwz9Mlb628rPFdsWxFf11tKK5COlA+3u1eGu6jP+Aeiag3mqM+0wDk
Y5HwuI2DeemNceJgUDW635HNddsmKE556CSkWMMt99Dl3zDzdS8n7RFyevtFHUCZysKp6ujiNQxC
GvXgyp4DvVks8arOz48i8Xt+KggeyOrvZRvmaPdwvIPWISBgbfwQzHB3HjVwERruKQU7HMsaTSYO
KepFml0khkN1QDJQmKmD7AHJ58eUasUpVTmacyLCT0UHv0mTqRJoJp9uRmh/dQMZLC9l2/j+e2Ju
onDfMP61v9rlPBOH3uy9+oLHwG5anhp+IsAOe3mFxZfH6YVSXKz5TTc2HZoPLNF+eNEUrREVdb2w
ehExkA1nF0xpmz7Bp17sbBrccWmnb7FMNbYu/PYIluv12JqTz6KrzrnMU19sDYU/MxIl7yfXxYix
rJWl8IqJqtbH01tHS5MVR6uqmVfatIiu5y8FskAUd8E1vWtjOD7rdk175v4S8rbSX0mYehBoHw2m
fl41Tia8y5xqhHdZQlAMfu3KeYUfO9aT8lqhetsz9eyN5tf8mzc7a4jsgXHy9FblSNjfJdZDoW0M
KCwm92wmtvSzzUqWRspcu+iqSmu3ahmFLzkyq9mBcVCuAloZJ9i5UnqNUTtRgNWI9apoo60bq7Ln
ilFOgmlbhnQhbpABKcET/3Oo0z0SVwYgc+D34Onxpb2I4EhltwiTsyyWQBkTzs0usjOMep/U4yqX
5Yt4dxxmh3afjEEeem284FVo61MRrTmIsVdvVA4UJFBbYBSIdj7UhxHuq3Rd0a8pSEoWAzExAHzS
KUpROx4//r0WCqRkzuFnLbUkLHGIC7BaL+NCSVsqIecx9HtJiXbvlFZNYV8S9pGXWiSVg4llXHIK
d7kKOqzWeXqlMxl9eUEGf6WCavxj5nNsPcsON6Rbx+CZ26T3f8DBIb6zCSjoLIVsV6ABhnMKyi7s
7GFpVAKzjxWpxy+4zGV9oIe22diI/3F06RrU2pHD5chPRnQNw4B8dvEHEQYS6Kz6UQU7ZWCSEKn0
esDY7Hc8foBxb7KYttZPgJFUWfm+o5cT0pWBURZ34ZcbIJNjOPsyvBg0t+ptH0onVeHgfyCm5gAi
N/BMEuUpHvEeaKtQxbT2yQw/PItPN/Gg8HoAJmxiM1gO8rV5tHm06CQQu2Rm00FSaJwOoosZnmMk
A1UywzOYe2ejaHHk9JIz2hCigPQAU/rQ6zM8a+nPunGHW3DC9a/2V1U0dyWV5rZ+PkVA+6xZLqaM
3JWBm1f0RctzJ5PeYNBPwvt8wJRGwZXo29InfPigDn42K9c9+hRtDvvqIn5pUXugepLjIqDuDHHa
yMuvgeU2+2YmnLEvhgOw0vMRJ2tLypQjzKYIGPsfSPxEWxW9ibsyv3/XlNNhzyPdh8jwPk9h38Qw
5B5FFk54qq1y+DgxzqPHJ5DAUCysXDlFqxz+91kDXG8pubXwzFMS+g0m80e7qHUZSOaenfczFdHN
mKYwuU5kpg5q3mTGgIEI9QuUXMQ8bfTrobvkBGL7lKgQ4FwesLigQNR+og2g6PyjwkFgS+K7UmdC
bUQkJJAeONgXIt9dWEbb/yeNpol3QbYivd0LGrt5g1n0+vNpASJAlhlxC5sy0rPkocPsNKn9xYu5
MLQ/pH5KDuXFmCHCFmiSVmRFbF41vWXKQYvgBenUnmO/TQ9nv95eaGyJMgJYp0H7EGJeUcmN9Nxa
TowzrEskUkdO45EqnoPpxtp2i4p1NjVgf2NBiqxT+xBC8G6s6Vk4XA1mhOI8+LADRApI0KQYYfJo
Qv176ASCq6H1vvPCFZa3jazRd1nGH/zgjtawzYaq5sO2h1bxeNOGrs7n2nY3etssFJ2zwsklMkyW
LlDLs+eP62rxSMnRec7L//7B9biZD8S5NLDMX7sDV2wi1miBcz2XmUun7xcIhm3SCK8HnuNtpOiU
3yycOQCK6TKK8bfp2zFUcmxV2ToX7bmh2ZI8tEJoVIkw/5c+u2YMjLpMY7O6CKKPpjOJ8wSIio4z
p8Ac0ZmjBQKOaRBIbQaGS9QpHFi9YUpWebH3I4lgDwqlkmAGLUXM0ZoE1U1POiQTre/Nfl/S7G2j
A/Xi+P20pLiq97u5wg8diZks5eIYAQi5TC4pvygOehd8el/fwE9BERjftapr5CNx1/44qBlnUzyO
tHXooms+lkZe50novvuzGNXr2sBaGZmkqoinx7cyBJKSbx9mKj16qasunisCKoO0Yu2UKgOwr4vT
6EbqIEvnbtNokYs2bgt6stcgOjhpW2XbSLklEuAx9AnReRR8b/eSmtP49HqLdtzw16J53PQ11Rsz
i5jwUNEyB/Iyb22S0ajEveG4ObGEG2Mbqn4uEchS+mmAZvpg3Lbd8Lkv6FvBqQD7RenhdCzgIIay
99kRPcN6ZvN74rkLvCGH7tV6GLHp3ZkebtEu7c7C1SOqIIkznY82vz3y8eojpVmQp5sikdZVPAjT
khX6lSPAhXGuH4+zVHK6w2DLueOZJijAr4mqfgNoznQh67P9Q2xqno0odIlM45aa23n1rGm06sJ3
unqHE0Rrav8ZnC4MqjmwnVKZx47+nxNqFuYGIdMNxzwNjM3kb76AfteSjeZWYHqinrwDsnAME6bz
MmkcIVgVDIJSJ8dRXlw8pamaArFg5N/c4g0gy2JXybVUT4D8AqBlnXid9SpbHUEr20QY3xf2ayP1
1D0pynvhfHXJVeD7ELfqv1zYUPEOc6q9BZzKvFlZI9SuOQjL5I3VEXQ8AHIf7yRtliEVIkNFMoND
nW6mAP4yNBbVuUmIP2pbwTvrnGwL0RWQWFGswlZgiuL7x0l0D94IaAItyMHpM1MUqFDlgLGBjzeI
IHf8shJrVlQmmM55Dm9YMswSq6A9cSz0+m+4U1SkiPGe+jbNv0+BZL44j0YE8i3Fqt+W8lFP+h7C
auXmqIzh2Khn0qlMpijoJJZLKPcdKoO2Yd2VIxb2Z28wgjiFYWilVVP2LzVIO++R3VtuEfmZSWVW
3Oc0v8xQ5N0/10FDG34dXgYv1B1qcDszIUibbymXuvKxepd5fq1EbEnUKMs4Y5W6MtlnGWmCQu0U
4Y7iiew+eKK9AYyUC80eojmLy23Ut1mWQZbsrNEv5fQIYyXOvwBEb1dpVj+N93wfMQ1NQLy+7CUy
T5N23iClBGfM+G5XnjJ49ZRo3JWSDxJlg+LfMLuXdpWonH0Yehh2FDMr60LuR7DncVxsYXENmhZs
IRyzv0QdubYhjguzPxQaqVAxRucZDjrw6uWt0FjcEEn0PXSvDp0L6zG1frRe7gVpnGMar0PoLGQK
Mk2BeXgUPypnOFlq1rNpBKJl7Nsmd90ix0GKJDfxeDW3x5S9rwHU0M/2Te3L5hiLKhkN5YPNb1h8
2RFy5wWo5sktItLQYiRHw1bF/2V3wnvz8w44DqGm3K9TdML3AHSgI09xdazmeLsaeJAT+wTzryc4
Pf3x9x67MPxexKv7D2qoCly702oWXtNXoVBMECLFX/nDGYdG4S4xTB8rzbU7K+tX31vPlvihAQCD
vOgnrgY7FbRvYVixWOgdso/by6DXLZ5AL2XShNfQXKyibu5wFz0DB7VAOnNu8kPGHNXg6WRsZcRC
VZSnTQx21B8jeDEDno8IjDZNGhUGgU1oECOf1NGt4hhYOc36n4OYMlfUVLL/lcL6n+15vFBMqEi7
SYOwBXOdQmuaIhkhqq1T5oOygSdtQT0GPZ2fmIAHAPtGnKqbzN85jcXy2QnQiSxjMrG8N2gvGexd
sRPsB+pIbqqe//J60J1pPpbrfBJLCQaNB2s3Jw9o0E1XG5Yuk/4iBhMNCkpEIcFqWWKSR8KMio5Z
pwLilQnFVug4JXBrGpsc4k/ulY4I2yn8ihQGbK0+QvvnLPo9BCEfqWkOC2PL4zjB6vjUv+45Fio7
+HWXzU8zMqVJDUrGVj6Z3RQyhg4Q6ByhXrFLw4BKBZfMrjf1G4JJJrjeyAMa0soWwDWFqUd0oyJ4
G787t+jqYJEl0+JQTWfOsP6ZfK7VJJpLdho3mHf/RHpCO8xV3i8Y7JwkXwhiCdcHVSR17MsEm750
iU2Yu8ycxN9XGDPyZLjyRJ//uwRtC4c8sUWlZMmzLdc3c45OmYLGMN/7MdAHf0kizN1abym41m7q
E/67EmRfA21JlGR7xYMLRE98oP2irEd/AJLQL8P1TSRIJpvp3zRSzOURPSRS2Prw4dBhW5Ez2LXe
iJ1wuXeYh8bmcs69TzwOoO3TULld7gckKkGKG3/BPHlanqTPkPA1MZy3uDXtUdiLsgPuTae4aLj2
2oA72ANj/YQNxH/2PhykJGbO0gq8C9W7JOjmL2wDOFdCNwZGGQkZQxAsu2jfCgd+AXz5ji0J8X62
iTEK9SH9jAnluHygKC82SfXvNwHJQ1/A8n/+00yzacLm8/SlVWEhrqUj4OSOWHow49bvmYP13bxu
/yteQ7QqWxnR6XIuJFAX6+zhFvWO/M2Uk56P7LKepEYqwi5U53MIXoRscel848yLOQCS0JshWNY1
Bc7g4FW+JewNLVe7u5p5vQYlChxX2E6W7nM39Pb7FXo2jFhV/NozC2yjuyWI6CPO5vY+RI8sycuQ
u9Rc6reKfuMHEqq3uf9L6NaWtywxat/u0mVvMWkCnF275YM7oYZeeSzDM77apz2sJI9c4YBxrMA/
ZLFDspq7Ly6LsqgKqjcNS+eFxNpiFmGEJfD72x406bI3tyjFtcwNOyPTvKq8i1nuDL4wF+QKTR9Z
T+9kdijI635EwFnfzKhu2wolSlF0esJush25vFd3uXPxXGn5dZlJ17pd9hEaheFIevohAVbc5EJY
35FJ0naJe4VDP+M2vaQkJfvj9936xBHbLnG0Uh9Wg5Ps7kjOhM0Za49A4Fwl0u64rUn8Bk3DYvq7
vtPr7pcFILi3P93n3rl6AKOQHIyMQSaev/mfIziThV0eOgg6p1zDLU8PEETfBuIoxrm+3FfrIm6p
AbDTOkSi0IIHoB6DcLXl1D2+kOjyRUd5NzasOFfgDEB0UJARzaBBNrMD1xylLvoFZk/6FUrqaxeX
7Ht8c87g+rNX4evi2YF/fhN+eEZcUtT5Z77YcHZPkMzsoizawNEzW4VkADuvBz9oqx2zD3ZcZAEG
tpp6EIPWd1z/ffBvUPerIl5mgtmkpbHb9loIskG+9+w69sNdW1bBP5tLJCM7cDozjhpgIjUfGo1s
u+epY/h7Ilr++Tl7C7L5k6h8EITRy+1GatzxOSgUV+VZeOMmahwolsfQC0cUMYdJMlcG8C4Tqz7F
rxUkyPAhsWijakJ8N9FDS3fAiWb3USp0+iCcskWh+x6b2TB6SW5omq1a5VECRwZ6+H6AVVvVaB6g
3RlkLWi2VEeI3UkVNlmJ34P87s0tCKYMI2JaimaiLilfBsr/j/k5oQZrZ45J68Wii44ClrrVzVu7
mFjtXqFmNMYhEE2mLiuGC7ZovbNxfKlT78nybuqD7IJRArGD73m1u7AcwW2UBdAOadL+jQTlM70l
6Wslk9sxCZQLXJmXS/QATW2XOln93CjYVqmEyqkhMrlgZ0Zx5xyjtcGqy2UMkrNZa6ZKZwWFo1ng
U2HtcwqWww+31yJlWdeChfsviml05xq+0138FgBxEW55YISVVAlY2mIynS6jm35Ws4AnWSyD13fa
JTKXRhgmmzwkElhdHP5EYt+ssjGhbiYDJVNsjpbWyvWyGut6ecznsVhTyjZctCbeFtB0Eb2A5pcr
lNoUBX/JRbkNc2x6HdLCvWHRYvX29dKjO9DPs55Cu9UHnTidH8EYGH9NWlfeNoVIYd7MjfJ+yS7h
JvwWjaq8bUoDLFLGk7Jy9T8a3ApwCjaR1U2rjqv/7mqszKrqXQwD/saFtv8VUFzAG0skLNHLHWiq
9IFudgUNBZfan8nQDSYLfM31UBise4qm5oowTQw8z4ljxk+KLT2o26aCkYJgwC43Pjy40gxpA+5R
LvriSfkAc9KBT3vGRVN8U8DnW4Z6xlTd6s6IRHJP+tYe95F1lmV99nLL+xx3sh5iI5IHukWxgy2e
FPpXYZkKPK/3rblu/QnUA6N7De7MSS3fLjn2PgD/+Fc5Kbc+qrhDOsp2SXcnfX8WyEa5gsbepqmP
abJhWVEG7Yt4alGBrdD1W63EDRVfOOSj1oxcJfDXeUv+7W+M/CmYfX4zMJ/G77WP2/cNR2LMxyos
vuZ+hfIg5v27vHqubonckfw7q1t4sLJX4txIZt2MdrJwkwpHeeUCOvtledaW5CVmjA6VEcJfqNAp
OxSIrFXUe0gN0DeFBmxf/KM1rMFHxH9n3tN1hX+nluOzMR7M4cmn89Dlita0+TkQHkveGqkcZioI
AXdzqWJHyK30yua76w0b/JtfSY5Wt3omGW1bZmcUbsz99HNKiTGEIK9NEWjxAiA5YH/TM2dekW8Y
ui52fz/o6YhsXQXvyqYwSbZQazYNn30Tiy6y0vcd/C+uYSuMd6qf5WhjTqD1K/NhOR19yW/eE0D6
ZquiUUv20RBD9uNu6JNZWcxxFzEVLzfYAsMhO6F3xudrRLS1cpT5l+TCanbKQPJQx37aQMdtbbiW
GEb4mNFrY+4lJB2+WyjqaFtzMyHCKICcXWevCpKfTrgVF+BrmrGI1MgDzjg3umdbyjdx7eHnp+c0
P6pPbGC4B4NDrcIUj3Fll1qMYPzH6jlGIWCi/0sQEWWD5D4lsxUxQsRmJBMI7j8cIfldIDMAXbsu
gbfgg3TCYr5z6gbUZ78uz7LgH5pVGTu1wMZhU0pKnmHKN/hPV8dIKvSyy0CjPbrN7H1xGfcCVmVE
9pRcQaGDisSmrwT+6Nem5yKzVUxbgnjyIH1XMyMPa4qLqXErTMqpRQjssLqFd1hdeTFV3ohNFf5L
LH53VXUMisdFl+b9y86r8eyLR3BlbND9dsd5fO9ksIJ0Ja6mgTSkTTeDxDahe35FgI8vDfGqzUYX
kTdPF1BlYongUv/GUwqPulCOGJq/KgBNWAi4rrkJeRy06xV1U/ZzK4vwsPlRjUeLs4esYM3zMNdT
M4hDs8f432czP5gz5xJsuG6IbVNdK97/GiWJg9bIGiCLL2KucAPZuMNmgh+Bmf6S28e4Oc+WJFR9
WzTZqpGlra1H15NkAqp8t/f/RbjRBVO2NBYIvNfUbiCCpErE6fL+K42uBj+W5411PxCC9d6ofGxj
eDT02kUqY6VIMUbbFEpwLsRaHinZVC/PNsNJQjNYehv3SZbxxi086g+U61wHHYoQIoOa5QbSH16C
5zlx8qrLx1Gf7gqL8K5oUsEKXs98aG/hglL04FOOP/XfEkPAv5SvojWXBusGvtUFWv0U6yfAQ7ru
mjmoc23LnnmLVYWFcAZrFwgZ+yqYh4NG3TbYY+MPXr1I2xv/tiIRpwQcGXYmnpQY74OLsniVzmoO
1WagueVzBquyy0bSicuk7S1Kd2QFsbg9KFYQ/q1YfMZscOvo4WvimjjByq0IoZURlSwYOj/DHDjC
Z7TdLOz4a4gnNdX0j0rzAPT/2URRqePp3eurexpya1ckijK4/lEIu3o1GrQ2PGKAt4qZmBrKQm2p
Y7uYXkjW6ufWN0yfIXPeL0XGVGzBJBE0m4VpLbb79xAHcL9kqOmQOzdLZsPGDDI6KiIrcHCqPwqa
E8ZOovZ4+Tm1Tr6tsK38fCY4YIYUonSqmOPZ6SXywwzYCPpKqLUdqy1hrVYz9zrKstYEaWmkyKOI
18dn7mf5JSUl4q3LIf3v+vcwcu+M4zoKau/FrrP3s/XUXTYbNDfChzeG3Z8tt2pI9qh8oobca207
2Z9r0iaaN9xo/LrM+5V9kVi1zUfUM3wBH5kCTBeJ7JbfAC48Q8/bhZYrnaBa+l0/aVQplh3KVtLc
MdNP5U1pOTijbhbCe/idw1SA3jeydFqxugMQwngmYeLNtyBthg/dkN/lPA9sb1Yl5YbUvdeuhkxv
nKTWhCkuVJjJai70oXkU6RZ+3gM3/bzZoVpS0K252r7GWcRCs85FlHiZHQErB8R4SVOsLSmVrPRg
SbgSnA0iuHBrGELE1nNtSQ2n5pZwTKVOFWjdSipMUYRkkUR3cD9mM3uBgWJenAbGQLum2BM7HLsZ
gZRd1MLSI54vxyeIofyfFMzDHcKOoNLZHJrXlgPWV8272mU+HBXqoPx2PSXJLCiJPb+PxGPyveIL
2FdKy0f0BZczgdUIS4xmrtRz6NQSzSFzRHSsAYsi/kOMZtm9FOohKVNEAQLg9PA7syja7EXtVN4l
IEPJ8HTxO9EMD51P7ONsAqircj9dvDiITUnYQctkn65Q7WwsYP+B699/l6mQndzmkrFo7UWzrqxw
yIGf7t/VBugHi/H6qkQrnJG6qC6Xd8ansUrwA4BMh1vB09lhJCe6NH0inBf0H5R3XcUZqD5KmBJi
qOSK470Jei4/UPU4jENEGPqYhYgRMmrz5WQ07O0zZB4gdr7Eq5+Saz72drBKxlv0euGK2I9FlZmw
3yPZ9gMfC4h+mwykdx9MMorKhy/Vgq3viOYfiK/LM9yp/J6K7w2/tSoAWFDHuWm+Vb5P4fEJJXTD
Ov3PJ9I9m13A2Ub4xjBiPvVR7kIfoD8RWL68OW07hJ6/1YxYMDaAH0WdGS04nvV1q6FGSx9mSu+i
jSCKp+N8WbCvsT/A8YWvGoLE9VFfZgzZIXFAhEfvF46IbCd4yFuSdvo8JWF4hPELaJ0f5ku07ukn
qp+gFC32gBKoAHgmOuSZR7eP5cJnMeaSq5ph4xtRAmCR38Gk1z5AVjU/Nz7exrMoFZMi2IRk5g9o
LiXeAQZxrbt8DXuJEOh/HSd1wcNptkiClU3BqSNDeb4UBDoAdyLlk9l1ZeF6ZNwlDdwjDBSuDaKW
dVkpwL2sf39EUsV3KlrYSKJFLMHuZTKABCRgHhTLX6LFxvfN1y9wxUw9+kafUVXg8rfOdnwISOxI
o+9awh2639ZdLpwvgz9b5ko8cHkcxFO7oAz7dHLpNS38z1LKYsZVr1KFudJEXKi563QgePX2xfxz
DN3jPybAWfIZ1iJBJArUNc4GxnRIRNpVUxOqTWc1yWMyFJ4qNN5q0tSHRlYXQ7aousSG9RHBfJlW
UQvCIP2UUB+hchhoAs2o9+D8eRrj2edAp3FO0/PP6P7YumSVKXT0aHvJpVpnguNh9Hi4M5e+fiGz
O+jtFGjBW9vw/74Tg/Q+wwTqoyVKvB+UtJ4FMLcNAthoRWgHBgdMbmqqBboN+ozTReUt2Ey3iW5s
v5arY7B57Fqlk7aX6qSCGOy8FXtq9OuTn+mPZHfAa/lw9kNGVXAm9tRsprn9O2SuHR9YuJyYPGKf
KC7eEC+iIaplVToFX5M6fY1cp++Z5B6s+yaJnuK2m3i3IlRynIxVlkiiJtoDr4wMCwsSC92y8EKk
TILa+k8CNYEJpvWJOmasUIhGUnZLvRQZtq6ZC9kah/g1xNzP2WdtoZaLLZVELI5Lgm3O94tYKvQK
1D7RdWi713lzBTrSokz4DskrMLOagfoIG0HoXOdNZlTJRcNKt7FsZ6yuBri/UoQ9OqPgL530jaa8
s2yzufj1mGwktq1PHqTXZkoQgS8pjXHE4VrAoXWVLAmuVKijLgeeg6GKSM9tnK8FDv9lilTpDKpz
jCgg8Bi023AVxshB+xFT5ONOESgQBYkT/+8kXwnvPdHeGVVP28H7ef8i5V67GSd5mCUukf9b0wG7
2XxVxApbBQxSZl2MEXEbU4oQQ8EbZzI6hGe9zDDJED0RPaqmFNgA9uxQCGtrdwj0Rebos0/DdGNy
dbubi5G5mSmLnGMqgTeDW+6jjz1zWzqo0zP5OUwS6mrQWsMWwFF0Pmg6EEbOB8vHq/uOs44CxgP8
B4Z647owuDxYrC9U5t2cS5LmebVQXSRk0nvcQLbcCkO5v4F0OjQ+dSZmWxHtp004txisWlysWXlE
2LIXssRtwmisuupZnMhfrTYty8d+XANXkattAWc9eG+1RTBFg+7N0ZkrUFIyJsKH6er/gYq0esOO
5NGq+glH4w5Jb/W8cC7M+PNxD4fQmyS+eHSVJ9vOpQZok20ZaJj1PrhCFIw++Rp7y4bHKkM9pY/f
QzYBiIQVoanNRIy5KRny9lTEOGPnBzjZnBsuR6LWC+1740gTQhIWWCczBC+jdbj2d5yS9ncneeSd
mJiOjFd0HMoKQl7d1+ORH+6UdkZhkjN/uruLiEFN/tcOQRsp9sRmC9ueMvcjFzRp9brwHVBn2l0B
YBtG5v8okopxFS6CIldP6MgPtSQeq3auvuh0aImXLMAkITjgWZ4fQ51YvdnnJ9N3zozO68natLif
ASyLqkkvkueWcgKXP+cb7FlbFklPIVpSwMFbzREp5ORL+xjV7Bal6bHisoM2qyeT4ggBgoBDGVSA
RTQ6Lxvzg8oZ3hK94qQzju5NYJ4MtsPSVf/IBd9N3vImBbeqUSUuaPJS2ns9/htPEk3X10L35tDc
XRAi2G2au7JP97z1QZdExa9w77OfCnJHTsqqRIQR6r5uEnSvsX2e0A70P4gV5tVhjvPNfA2SGb7m
JA7F0lZRqpqIuDQ8JM7C+OOF6VbrZPC1VDdbuAajuegcvMHw38jYmcyyo2oBj7shTK+ZgZeruhOC
msq/cofpr1bexjEPXzf7AM0uvD8/+oIRdDSTkJCuXOAYT1k7BCoD2tUeQ8sf63Q1lGqwkZ3jlzYC
Nv5TKw6NVGGtllXAEdxbTYslwhwvI4Ue6u7dSxDnDTqKUVENyDZ0n+rAtny9mBq4PXfXjN3vHIHV
3i2aVj6K05TmTPTJtwACNXXXCUGW8lT3DKme8Hbg6UHjdkQg7pwJDlp6r6ctqS8s2poco6yWZO2B
sv5y+CvScgYvMMXTUlZJkz2FFVwr2hnJ0c5GDIOVR99uT0WzRKshdJiSPkgNE+PtVO5da4UKT1Yp
gvJjCb7W7qlPYmDchlwXEgqVNXrrzJRVFBfNQqjhXHUcP3WX0OkEugEm3vqbPUrbBa0uVAWbtFXo
f8FFUyXZ5I6d29J4zPYqqmSgohBN77jXMp120kpI0H2fB7j0Nwxgur1+tM9hRsx97W5AfFoBCqxn
pcyyQLnMBe08LRHDGxnqxjjzy4UJxctofBAjnThhIz0lm0W+PnCUXzy1XeZijIGxAYkOdEGKlYGE
TbZGahfYviuFI5vxunyqNMBQNHDgTlLJpUaiOxpIGMNgeD4CGhmaB9XiiRa0TgFTwjdMaAGscr68
/z5BQ598j4904aZQvxbrIP1/8CcztE7ny9Wo/+5uYdICaY9VJyUO6vgxhJQGgbDa00jCXGz2mJXQ
mhFsB/FItKAqlr7/JeBU3Rtvw+naU63ECfm71U7sfdnoHUCkQxv18Z2CHHU0dFiDF0iZZ87RQWVn
x8PzrxM5UaMsleybNj28NS5D5HdDzxr88fp2XWVQVnh1w9pVXnBH7Dsb4JdV14nx+tQbh+lGbNep
YjqJ/Xybt7ay7tYPyhB9uDrGJce7jhkN75Ti9y0VMyqIHFNyyPnavnTRj/6KvHg/XauUphSvLGTL
k5+95z+d3K86GVfwt+jJK/BBFA4Hc1epNn03QyWUjApHgTizfGNnt4LW27YB6fpGEzT3+SiqtSDQ
Ss28V6UXX6Orgm7m8k+q4BWR/ODgFiEyr+jP6ncBL+16SRITffrTzlxoi4P23VAZ3xY7JpaQ/pf1
VkQyTqeW9SrjY24hBYLqBDyvblP5/KLWkHqe7sgkFKLeB2vMUk9kHmiaFSt1DnXqvw9ht9JN9Dvy
F7+Tj2x3k66ISUEAJIYq5MeFJqtSy3V7pySpNRisQp0a4+yYrQr90xlBqTq7hKIiEJC/RPTIF2S3
o0jJLWMD7oT/qxGDukfYJRPYWNsqPs6eWr08mVVE7gp0EX6ItsbY5LYy4psHnEZmarNxJJ5HgF/O
m4aEaJL/drj7EkxJ0S4LF/LcQfFBRFJ/L7oDS0fwBYzPKUkahlyAr5nhKbcjTevQJIgk16s9ZTWm
jgqhllAJjiw4BCXuf36SgMQpLX8wHaA48mbBYfo1832PGtHwV5TlDt2yOjdxJB1kx2KFGMWLS+ba
GGHbmGYTyIW+3O2JgP98/GK+6o98cBjXdKvGg4j/0qx5lUKZVqobYZdysTu+anwo87q93SgsOkHO
J2Q+bUd9KBNY6gCgQZjt1mYAEX2IsTHYIa0fCLoYpJLZ/zOTrdS0Xl9AQ99HEHQTIcWfjSx2n6Dk
QnfyEPSkBgGs+6iSPxBZeVwWcRYXvpVkU8OmgIbqp+lDZ+1X7zuedgHggPYxTab3KPDBjPm5SAyM
LNE7oI4ImFoHkRE1RtN5sEULGG1g/b1IVcqneQ+4dS9rYlqpWabp7GmS0nERbqpxbGTeV9GQMVVw
IX+6yBr5SswDkVJJsfrGpv0tOtiVU8S/NxfarReHJ3oeOVaBcBz5ditV+DNZmQBrvKyO9PEpzS/l
wbaJH1IxPZ/IK/dR8XMiZQj0u5LaSsmqQDAMwGdtXgbH7on/Ux1UmVBVTJAWWKyG+Ox6GMJhHCqF
an+ILBt/gtHOTRzX9BdgHkLxE/D84rRzZMj9zYPibjghAUM+NuzGsaN45J5KnjInAdWOiDoDLOin
X0tXr6pi6cpypG9dKr4qaFUy3uhjHCKd0hbo59lmqvu8EYmDwO6i2R8XJ6wVWEH/u1d45GI2pz7K
B9F9aRfiyKAX2dUqolisJDMIcfjuce2pZJwT2a2C9xg6BjnqPll2JYjgK7x19PuDy2qwEw262jp5
pGZwRrMpPeVTozaxInkZ+/eTCJ3W9CPX5UkQ0Xqvn+ae9wFF6tOCR89KTS9FpuuOEDtTmyLY47g1
XKCW8APJFLQboAfu8F3UPZExenAPHoFX/IE45iYb18xQQmmnwLdFPB59XUkAfIDAn1uO7GOYizXH
wgFfzYjucDee9xbOh2gwp+p4+U85qXKi6ctni0ANr4lPzsQ5uwuUV8cVlBsvZd+Go7nTS6rjg1zt
AgaTltudmDNwDmtZt1EyQJQb9/fQdVmZAUNmhzS+Gr3lZi4/rCHAmCXZOOfRDecXZDdm9JIB2FXC
8lfxXmiCoY7Ayl2H9szYrxPSS1o7hACeDy0mLAU8HLdDjeVRxpQv80N0IVWhg4w1b19ABBavnGOj
Hd34gsuOvDfareSSIY5TG38wwoIzOktq3b5UOEd4tLZyh9j5yPGzgLa5eOJ44hE9xEbeVuuVOmD4
JTlFFVkyva1WNSmi+t3KoHGYQ3zRVKoAS6mvDOxdxEjl8TuqPp7jwEaXRatvkeQO1EJrtPsSRaE3
xLbqEb/D2bEDRDqNKyaGiFJUT6phAxowUcyouzPk9SgRYPO+J8HPiss5aOGHi4oiBtu03y7urvM4
L/8V2Gfi0AYbnt+OQRl/dfTD7VCUvefQDgvuePLi1Ain4p9wehhNhqYT0TzEBz8998a0uz9/ZFkN
CL/sJJWv0BQL3nvl9PwVXcbDpe7Q0bcfvkbhldy0+ApXCgS2iQLR30chHN/zqeY9DfMwdbO6tJRN
iT9ZXUwLXNxv2Q/Q0Ih64th5sDv5dh+D36i6Dg2oZ7NLPj6tivOvMff9vHnGvseeGgHBPJZ3jECZ
I+/BjqJl2aBZGA8euc3BmfFcG0oytAJFr6MAhSssantBxacifQyeu/CDV982q0kWyRcow3BHz/tH
q+FhuZryOPDM+pXNgCxAjZYj5dzwU20lrjESpyY3QYlt1TNZxmoiErKa0TQFF/kyqeiMoqr5Cyip
ByMBO70rUnFftxQdPK5/IoqLNRD4vC/RfKUvhJzMcrJZ3vdxiEEQm2tDg/xS3KweGuS73MFdkDWV
HPa0u6orY1MQMQO1RWV34IpT4KH0ifRs8tdsbKkvSS/IIMkwnyfRBUiyH4jFV6l1cFrimMlprJ8u
xxs0LkpAGgMctFMsx+8Qsn6hx1IeaTgPVV/fqmmPOKMG6cU155RWhkhzohFCBVJOpsNOYn+B0fBS
apOibh0rUEr7ZvXtJuzecmgATcKKheJlQkm5mpK6kGBny/gmKo1iu+c3tqP0gR1mPIv5+DICpHUT
iR/MASdX9kmqjJoHI8IBByoGyMcdGegWPeqN8/AdzOWsjDQHXpepylMYhGslehMJ7CEdme/6Zfo4
tOxeERiuRJi3kTq5WS/B33HoESAHka2nTNf1+j7s7N/5piiTQqkfwmmYiRE9wslMMTqy4o30USTe
RgsO17cKQL60d5Ph0PtaoBMxfCAh8C6VNmTBm0c6SkQjcgEUEPsgtS1B8dn5tqlJoYqgQLEVNS0+
IxLHok5swSGAJLhMWREh7EoWBO6qpZo81jX+Np8LlSbqRiVM4xlvagKXVrJB2KyzxblK9utLV+ol
/sztEkLrKnkuslsQ48/1MFvrgFbNi33GdmOZoAx5Rd30EtfEXyn215TgFbNhKQ2YO8awXPKixD57
19teWeIngYq5BbzZuiQMXlQTHk/D1rq3claXeSRJ3P6hcyuoddbdleu2DofyslmUQy77r5sbvDcF
jvlGP51OV0s+VCaUp4xzYCqkBWGLLzyMWUDGwe+6tdTN9jCMkWLlIEJ+4O6l3FI275Wyod3AeUDb
jDG4nvuWvkViLvlHRRH0xoaLzSnnc0lhZtfC8dODvuAN99eMQfjqhxqrcUbjoYpXkgUCRxeCFwoq
JXTQkqO1N6g9c3PrRtGVO3kngpeGp5i0jWu8ASXQNV0yqEJBldBw35VBmEJ+EB3KU4DLtkEXGKOz
ZrZmSJ6kB9cG1TWuOezGygbGf2av2uASmeYFkZzblPsvmnPC0l4yIIpnUjhYnZRjh34PwDAvgHvu
goCnD4MbDuKqae/V79tmE3e/e4A0NP2EaCHTZOPgdonPJjKJ8EfhD/KIDIJD07uG5Pj/pYsz+kQy
VHiUiLjAgDcW7jSmltjV983cNQViVXFotbs/NkQVyW33+TvkP80HXFTZVGzOCr7iBX2bQJQXvG5k
6cm0ycnjh0h1X40f6GBwVnXbXUaHuDVPLUTnk/JdYX/vn3tqi3CZdODN16wUMExLQdtHCT6B3QmX
7Wd1TyQRTuQzD8xwkPjmQgrSBHKYkNz3P3UeyERGQmUUQ6MW6iLReM5ayHa02fq8ArUydS6KGiH9
s1oMkbuOK/ywHdq8eQmeZ7+UAVVXuhy5f78fUU0MzQXvyRIdLDSbhERerndY8JtATGhKl+NU+fTU
ZLYLr67VT+coezQEFrIj8eCqqSXMtA6LODpaD4M8GnXu2uhTEI3pSRtAzXpxwm8Ye0kRMX8Bs/I2
FUnzz3eHwbzF8cuMz7Ubap+8G+h2wy9bGU9iDxgEwzsDrIEB2Hmefk68tLvvJqu3DR9mc+RnD9gL
wkI9MZ83VniDSQMuS0dKeoQsWjpY3SHvk89VUMUniU3qHVNpJxg7oP8QAl9pZPHjHgypbMnJ13IU
pQs4MlOxu270meIMJTzZr4+UVlhlQNXJxPF4EjfFGAjSI8xEXiAKBz3mdx8+GwKluoKpQ1PtAMDm
NsLj2ZXmYXDyZtdpyZ01RkXVU+xhnjCGkjQaP0qi/EHUlh2R1rUZsWEdZwdax9L/K6jRP5pawwFu
OFyubCTRF2QG1wJjXCtQ4Na4ydPAVhjIbuogU0sUOPOTenoNbY3kuZ2zkkYOy3Yi2Yq06o7+OxGS
RUESd4kri08z731ARBbwJduHLUTDgNkSoJmVTY5JWjKBgz6u0FSdIJW1IDAj24vFuoIY2Cj/vQUx
2QmO8KENupYU3p4v/9KiFBto/j/iBA5oqbHg2FrUsa6omekBAl59YVyjY/UxB11BGDqpJ3zF1RD5
DH9QZnDgOASngshUqbhITuKGuZzz1mWA1B4afPIq9oQJF63Z6G2cteSDy6+W9jDSlaO9uN7q1KAw
+TYzyXNBHuHDMDRnqt3OjJpX6pbVDaeJIADlDZ6qB6C6u604lxbtvcaeymHtvb22eXdES+ZLgIaN
DWXvoUm4id8DXmyTzk/AYOmCSsnEyO8ctHhsSSuSZywEZteoNqvdqvKVqIN7lFGwUizt7Rs+HMbG
d4z1VbR2IuEAlxZtmPdqjL2PXoK9gOAb6APhJVImYQ71wQRMnRKIdkhICnD5cbKNXlUrTJpnMAt0
5YfOrmA2VY6SbaWDlReQPcyLvcGacXblExSR1EdSEyktcYVEGBscjpEiLEhjdFRiIp5ISQcxVnYd
TmJcbfp55mnFAEXbi8H1dxYAqz9koR2gxH9EDBN8LhceyvqwEe8WZcRhvokMMGwOP1qcLopqyPr+
wTIRsUWaxNxiS6txa2xV5lbOiUz82ZF+Cf7euPKlIsNZNijaWbg3A83jZUlfPce9vdOSBdQ+RKJ1
s71EUaOavsUJxuZzHH5fRjNeR6UU1x5xwugmtEpihYtA/OK1Pkm91fWJ2Dx+3SIQkpNUy1NmofYS
mAiz19HSR3kF5rIuMO3urlDlcjZIKYRvkYXjKQcyjoUoS+hcfg6dPYnIbPPYXseOZs8ECOhyOiiG
XYKeG0S34IZmwybRDIblmE6Kq60mjT6jt+WywbXMz5UjBrz61FK7ik6pNV4AZZoWdb6QE8O7eB/i
la9HAclD9Vx3O2UdHLgfqCLt9WN6CCRySPrM4PCaWxcvU72LO2RfMdOEh3fb7aYCBbVmy4UJaEeI
19OjOS5MW59h2I8w95Ct9FDsRLiwz37I52kFouRLAuEmIr9++AkQ00Puqc6hZwCSwGfRspLE2FT5
vDmzzKJtizmC+mHBDbOquH18E1EkViP/pM1r/sJb0zaxCgN5e8ZEg3DSnXrimaNTn5X8+FfqkmUu
G7tBdkDeTs4KH+uIVYPPLQcPumlAs9xw9VYPuHJoQTPSdJX9LHw0ChDx47ScpRluZFTHszNglmrO
2y1zD1Pk2FyW8KeQvX8KSfSAMy14s954L1ZFNvycEKLhY8UebMyTjtDSvKTBNFlbNWxp8TMDz/ac
3SAJC3ecB1Ypj2E5sAOzMqkSdPVcQ40DmvLNI3vgtWQHnj1oN10Rh3kYTkGEVgxM/HboQWu/lDom
QK6UsUQYaaNEK/F/sTHuLvXkF3YZm+26nkzFHs8iV2W5Su9pHWcITHxUIAnnAehVPDmNc7StKVNo
a7gIAg4RwIJD4T2NMHqMvt3lPBUyeYDgduoYtq6XSeIY9gro2tSDgz52kJWVdg3Lh4nuFZGUi/UW
FOD7VgagCdAKe5gJLVLuqB4a9pojYn0Q8t85kvoC167dt+3tbj1ugeEssjneq4oclxXGy65smkCX
k8xIz5KSyAv6KrtyI18Q634YTyl59bZ8LLffT6No6iar+PKxf5u2x9m3WlhAKyIwOSVvlsu2CB9n
yJv33p3/A5Z90demm1RicSCkFlfqkYqE30nV7dXphLXYt2kujrcgxUoWt24FWMkPZwyrZUfdS/Mb
vWOVQStL3zH/36y3UjNFOu2w4/9MhHCO4gATWif6Enu9rlTBRSDW3xyTPV1Krlk0TEpVnEruiwg1
1rGOgzexoueM30UEtvpZPNe2uT37+F+F9MsfkRIwTfot3uK0YvtwSSeG1hD4eDVlY59KfdYTeee3
8VwES/Dmo0xfLRbDyrvj1g8a8MvgK17hUPkUL5PkqASrHMLqBsbEDv2e55uypSJBJJ9ws2En9T6Z
xEItrNvfoRjnZA+avXzMTnIeZgcg1eRZTicgCgdcM83U/jYOqM37BiYzzwpsaAlE0rygZAlywhPi
eqjs3pn3VvOumQA8ikWrC5AiK/MHhKYGVuRhB5jg6SH009c4COgxgyJlHldqZL7/bqzDamLOg0iU
xsReSGmHSW7IWJPkSyE8nSrGv+guky9cTF65KQcN0Oh8AKCIvUnehl5ZcLopJ6r6doikqmBzW0GY
nJBibbu7rNCeSyGcd6v8MYAILdgg4B6o4SF5eU6Cv/YYnHW0Z3kxavZjqZA5zOJw4AGJ1PW49yD2
+DqRVFlvmRqnjav+LuKETHkeH7qRnBeYRorAK2TLDEdbRwbV6RDBiyESfgVJnVyoI96RQgPbWCWO
+i3v2Sz45fdoiZ751dZkN5pjRvQsErU189aNqdADqOaLHKd8SbrCNUPD/NuEDlpHZuYRPX9pGOr1
eq9VOGvufdvOSvx6hgKkK53lppPoWJqDCidQH2Kj8SnpgXcWflvBS4/8pqH4Y7JOFlvbjuJ9igkm
LFK6mjZ1cuv1wFM4nAYJMEee+DxmDeKpPx7xUjHUId0rlcHjsiUT+f1atCPn+ZGRWwtH1qrAMk9K
+TxmoElWSZdQoh4AufQgxo9ifbgs+SuU0/0PhFyNNzlapiijcyW4158JluaHQZuTIyj2G2Xo2Ig7
ZqG7iD1DvWMmdBEvD9B1LrlV/K63nnx8VsiJMx/Qqmh8IloHH2z4BytSr95UUkM1jM8e09YpMEwu
ef3kUWRg7Moq41Ypwt4d/LgXMmybontJMD4zlf74swjxyCZHy1aSTdhiiHuci5Cg7qy9W4ivVEYo
WKiavq35KpfgmJpvSLy0uVrcVs+qcvmqFLhz9f8mxxt+f/z65k3XHgu7X55lI3lrQFr2u3wTG6M2
X+dnSgSPcjxdCtDRdY9b7N5EzoSgtdZSkRMVcrOnqPFTBkwL4bgH2CEBreXrOB35P+x+X0nUsC2x
5gLf7hTMnPJNVNhH/3cZ3hvcyVdme4atBm9YH+EC3Vybc3pqayW8ms5v5OXVJyn2fpz1cZ+9D/w5
Hp2Dhlw/mWYWV3VPp6hyP34E6bOhFZ/Z52vTH6ykZJ3jnJ0hx9jnTfKXeO/4KpBSN1UwsjMYTmZd
WTAJGLCZSt44WBGxd+f/ZihMbfmiDeB5mDCqwq6ShQgWmqNcvT04nR5+xKGFOqeCgtLuwYE5w5ZR
d9yIv6vnpBWF93HUjrNUpBGACbn2qEUFGAAsA8HX09du70lN+YthZRHuV7nO3VsXAd9Ds5DyvuGf
seEmCI8g6mtZm/XxJU6EeLj4chaM0t0ph5YzCcjCUMwOgRYYfESwlExWiTijozd4BGy5Z+lYL/rV
1BXEaVZ9jYdL0IwVCh5i38MKGRzp9AcCw8/ewvANuqFweUyhppDjpZA4zAiQgXqqf0kaYCdYiH4l
jYVXP7MBZBq+HfY5FrZpjcRWX9+e3emrk6dfc/MQdaAQGyXR4PDIiQdfpDAbRAfMUX+pLh2DTc7p
gLMDj+Pdy7RILHhf87ls+F2EeK4+wxO20elyjDVR/+MY43P3mvEKJNtV5Yptmv7yDdLPU2ShaFUk
lCQbEuU9rjZeOI5o7cPdTBT99eDW5PpKQW4FcfSP3Jt937v+mH61jAbWe7dQrG1ZTZH6cFlN957z
cvcOGX0LzvfzaoSzU4065gKu/LvY5DNhv6A484dBrz0DxQFJ6HC1za1CSS1OieT8oCeB9BHbbr37
H/7AQJV0EF9lp1V5OUGEpSOGEsJXHiEisqegkzdejKr6JZiXHjfCtft2uArJg5joMXAXlcCINQdw
sNWTBse5zgYC78rMq1KmtQqGShA9L0BlEoSLU0CVFzJOSlNIgxyg0um4qc0OyEKS2tsJEhriyuhJ
2EzHMFPg2iEAsZX0H3yxvshOuLS48UqqpvWWltZ/QCKmfr6g6vmu3ZRowYl7exrpuNeh+RXE1C9h
NNGcGORJC6FV8V0CSvGdhKfvQQhRUHMcuCllHR5yGE6GqcYNQCk0PUB+qnbv755zOkwinT0T1bBm
tkiibzR5F1e1YFweszG1J6NAwudzNYqnHxbeND2KYV/0+3EYpmz2ayXF8ixShejnS94NN6ek9Snc
4sXQ5QhTxA7jO4M40+4mUCCtXe1F5pkR41S+kvLjL9BKs0GGyx6xMUD+gD+XPwu2S1n0u4h7PmHB
CrhO0Xz2UbCSGQCON4G73GKc5bCXa2Bz3ufnRKIchFKTSHotDcHBE6MTtv19XzVyxNGJBB8a5svO
NLRVtqLPgGN05O/JPo2tis4+VE6hSBY6rycROKJSBSjqBtSjwNIDJQul4xuaEuD2TqSEjM8Ygh0u
rZE5gJTCI+5nBjopKK5xgFpFF1Lw8F41UvE2VQesWaGfNUcczpCHvZy01aH6n3minQSXmi6AUq1i
Rh4XKnwENyX6lVIVQWcVnIV3cRKSiP1AqVnQAIx2MQT5/CtIPdqnpEA7yB1vXtmMpkeqNtB+1Pj+
sWlmqWgP4Ly/pJPCxREUYpkeAUK+0tbqJr6h/ef8om8Ug0KZcTolD37s4uESEP1ZbYDgNZ0iGZfl
Qq+vcKU4iHY37QCSYQER4WEOeNsK/6PUldtX87uF5yFp00yQftwd+FG4RQddRdS8oVKK0+ABJCPL
QwlaqFQDfQhGhcBaC8kRG5MveotaXcnoxsjDG2DED7DT87tsghdBEbtD4SVsHJf3kZ7pHAm+ySmV
U2E+YDs3dLboPOQVUIXuec/OYkhADx2Chga9gft+vdFsURXkLGHovvchVKiQv4UMSrWhDD63Ll9a
Bm6vutag7YXGS2mFnyt8VO/ouM5MGMTEn42n3vUBtA4zOi7gBKbSB2HwI545XnJh4kSacBuOq6y5
P/fjSzj73rr+59Ov+uAkyXmZl7aaeiC2zZwSodewKil7d+prnSHomNTOmXcECTXclBqeZmDx3aXm
cJO/5yqJwF0+z8bi5FRmZTlbGvWY66swA6Y+ubexizkZyRubuzVdqCV3/Q4/hbjF1C/nh26K310N
Xjq1v7pkKm96FABYk7WIdOjaN34eypnxz3U+Dvcfy9axbE6jqzRxnWX3f27GPYr1q8o/JqcVgbHz
DBlGezMfReW3NrmNmM+9eI9MDk7ZBiAx7sD0iWCOW0oeA00EripmXivXeMSx5AYLpmvIU2sAbHeN
3vw1y7+ZACR3hEXjEBpFx6LvJA3+jqRhESHW2nxWh6YOquPAk88zWZKlBTkKsLPImJi4V2bgAl1X
cpehiSRBYjgBvcOCYJEjWGLyCfqrj4VwnYDNxgCB2JGi10S3P9nyvzGKp9nwzmDLTAZobV5MbKS3
uyDGlbJiRjgkqCUBI77TnyeivWPMtMzvzMXj9I7+2I/CzSGWI3XBcYUNNQf9EvgTaadaFm6XF0+2
sg4IlLOT5f/fgHGdLzYfEaYP6TiI51CIAyWTAMr+p7PA9XRQYIlStgsCPxl0r2c8IjuuIRH3XPyi
68XXx4PSyWmwPZPlCrWzhPiR5IW+tH9jaL5cO4mUCfCxLDTvMJKVCzoiTVsdCa+gK3R2PjTEqFXe
HBCK66n0uLlYvO+A/PuiYtIiaipalg5fcFhy9GKe27e1dbR4/g/Dt/ED8TFAIYO5brh9SSHf6RIi
iYf4gYfhyf3CefNpGQEVdl7gK2Zo3AxQJ27HUwm7xbHgpPlibGA/MVp1smX9kwD7KofnIiUNjXPm
rppKQgvz3NESXBbjp712jF9I7tCTPr5FTy/RlwVYyU4kDICrQ9Qons11jj1ZKNl1n/rCYGkevyA/
Ap2vjtVUN/rEolzhzLc0VD9BIF+XuUg8lzWERdj9zo5TorXJswJMLYJ2LYKNHP4mxUxBQNVtos//
oaWoafpdk8S63dMSLa7bTSjNXknTEfTvY8mki+00Vlq2sQAMo/vOnd5fudtRPVjSOkXXRtIW+3ei
oUY01nA6eLrgNLv7P/mt3t8P+zIbzqvQZcnX7RjJVLJUWjss5ZK5a6JS8Fzan7zpdu1ao21ivlD4
LVBeaxyWSrNVUnOWofADzux1Xhob2Vbps4UdU3ZTmb8ouCvoZRbrAn/39hFxo8hc6hhy1RxGKo+X
oi0cnHQgtGctEEc2SHaLmKxE5G+QZoV/ZQbdsYzldF+el8nRzeQOp+fi0P2/AoqL8rvGibTJmjT8
x3OJEn1OLpwEsTsU+Vu5UDTpZ8VL9wWLjrSHdHwh3Y74S3EjzsKboBhQRmI7kqinhVvvfx7U9CgD
2Y8aKzF4eLxZMkxZgEFfXNSlE/Wi+5QTy/TMAtDBzHgOl8LqWyWBCK6oWyvKzn+4H7VJmw4l9y5u
LJmddxeJbxvZlusabn9esRd8oIvW1gGxxE4BkilePimam+AbPQ85oF60MnsZa7Erop8bZGsSei/X
MPILujth9U6yIhCLuLVhjJY9em9AlkvUWePRhxJJtPC7WARY3Yi+H0sWBH/vhONGJGr9xxgXsEQX
6vm1ulor9jMJSaAwEssi/lhOp1J/GfspE3O2Kp0p5DitR5UnCI3ngXNt9fSqZHEBlTfQiD1J3/xu
ZeiavA59ZqeWHGFjyJ+s/8dig0fcR+Zea/g9vqUoyxcQvTA5zFXe/3rlhJXFaifEaFKO4+i8eA6l
2ELssRTx9BeQOx+IXbPyIMtjfLqkGC/g3q16PmQ1muccZufqu+W3k3+CxEh6VjsJQfv3HNDQtdO/
PtTzb8FTV8HpzK+3RGXiFsL5ltoSuCrpSof6j8xhstKK2Blbf7h5nKjcTTjPAu4UGUGJD8huBxj8
Lv4+blcorXTNc3RLatXEEbSlZagKO4DNv9DEzbRfusfVi1+XecpR/yE7YnpGI8rRL8+jY5ocFbnV
X5smK80goa+H7sbbZjqkt/lbitSMKhj2CvIu/gYAVK1ftr4KHpTmbfOy0ntik7LHjbltENtREThO
8bLt2WZa3P5XjcymFtEhskkXfdPZ/CXOVI0fYmZnItTCmYR2VIoehBJsepnONnI/q+QT5w2kLplI
4N71NyDPs2wZlWgZY9xkrejWj+/V58B6mv24ZZUXz4gd/w273BUm+5U7UBc8ZigwB1bmTGLH1IBx
8zrnvYhI2qLzn1Qkf8o0tqEwo2DRy6CEflhzsZt+58OnECMS8yNbXFVV5RcFYFk1YribxSTu2tOm
2ienr1Hc95D4wa8TqJgXg1XTWRac/5LBceQ2QmGAmALHTb3MrDvIMD4twGMXOfAHIBgRMChjNIsO
JPdDFQQs/PccWtDYI+aGFvfW4iJ4/nmUahFZLVyRlhVBaUoiIHqG28mZSHeGbQlbLQG+Nat+vbIS
UeqMH4t4GyBrV7z+ycZJTtVFhyWyKOjn8vHQa8Nn7QmvIAk5uGKCGYVKTcGJ68azE7jgR/TV75Gv
r4D5nURSohUJGIF73DaBcnqsrLYMFeIyFATti8Q+vTarNeyrT6nVWJcuHRuzk9fEnPPi3ag4SaVp
TVj+zu9pHoweFLmc47+U81OZwfsUYSC1YQnLwTCYCsyjLq/lU718296YwKatx/YLpyeavMvZloGH
AEdQzt8GwwL1o9HqwT9HLGNk8kRreRW10t6m50aBGg6qHbLY91D1pb1k/zAhIHm/XHqLJ+4GNdXz
OOOHmef5tqZEWyQYOAgzU3fmbYPIpU3YDW5oZzRksR6FLw1MgY6N0uRxF2r5LUiW02Btb3o4cvZP
rjj/UFe4Zc/6uFFpa7P4H8K82OeRTZkfnynaWI7GiyJqg12zCyx8rSg1xHT7pwq85Zj+G6yxgY6p
LisnEq8YGwgG1cj9g9MN8Z9Nr00J9qJ/bUp15LApU5o0bCs0baUjJogutXMPA2xXUwM/FcbPWmdW
MHViPOV1Vv9QQd6JmtE9efeAR6L6dvihKUHRXfJQy+vJTveU+TUnRGA3avClnLPnydTykLhMhQ6c
GefSMGNY95YkPLo4E+K4Afd339KD9dAiJrxn2ihRak0YWCu4ZPVMnPXAvlpg5o1ImaSJI68/JX53
LXFb+7KyZGBqTCnah44yS4v2L/ibbccKIXTVgCRJUKNKo3ZyLS2MPj5c25rx8/aNpG0C5X1a6TPS
/RO700JqK/GQ2vJcv0pPqZG1FBEGADktjIgkNiJ1C48rhm7ucmcroghrIRb8cbO4eNo2fnZBSRhv
0BNubTIzsLQwHXQtUQPn31ZHT2m4IiQlZBlbpa3qC5M0mJRxcxjDqyUF1fyyuA/MUMC1A/nV0gJl
tiRALFpqxU/8Kz/Ce3/7I7H6aJm1UYBgbYeu/thLL9cgdo0JMhOaOBuYHaLwrfsdxSKewRpYz7If
lueY9o0jExB3C7NCAtnv/vGYKrzopjPZxE3I/7Bc4i45FFfkO4LzBFTXEHAWNNqAbgYko7Vzel9j
Ybr7xp9WYzpEeOFtueuePDnL4K7WxuJ3Wdnx0EMIVAApk6+PQPFny9/tOxosJrzNDgj81VZlA5u2
2QxSi900999do0K+5LAWSbaurarrlev1ahums2BwTb/kuoYhgHJZzQRnyQVhorj54dhb9Zyzv9UC
bDi7ctVj5Z2UFMpB2BP779uMBaADjzZLg3cM15MR+c3chE+fFmmlv/yTJRvnY/tj/UrsfFFvDO+w
dJzaiOWrRW3C/1AjL5boe1ZLQ/EBUSh4dmX0IbBG7CbscPMri/DjkR16arO4M03fOGNXJlqIvNZU
lrGt8ahIGwMi6K1PqI3zI29rAYXqLwX1dmKwqoM6dHl6xxsxHzdKo9UqA5b7vZHpRATQm9Onaydg
F8p3irdXuGP/iKCxKEEtFElpNicKx2p6yq2Nhy2eKRr60pla1tYgjSBIAS5K7hFW1lmzH0PeZ0Xs
XKdVLcgQQMaWfauPS1p/kgA4vy8iOJZ8G0EM4ZRBGm6eu8yhDN0gMpOLpmjswfkSxlQdIXJ2LpQ/
9qZTIYm8MVWMumRVzkNR6wk8MkKUUBuKG7IXiKR1aTKGFMK4Bnq2ZqHa6w9qUA2NTac4YDvdBHLr
nQO+a6fuvm3eAe/v6W4jXm3zfmlABxnoRpUkZiPurjQKfWrE39QqiHZQhtmpn15KJ23aSwMxn1JF
mJFNXYvShKeoqLl/mCT8Itpw7OtzOrJbHYYMmi1b6fq3vyGXzg+IZkxziUDWrYa7OUBLuJ81JVHI
fo7g9vSPLNO8VNfccVoxqwgI76ygJr2synh2KDQ39la4EIy5Ds9zLDppNqXoFhV+zQF7gK/s/tdT
BvTarsWYwkEz0Gy/rVoiBGl7VfaGpl+qDtDf/3SPYutbH+c8oEkCc6m5ar9kcVkP6E2Kg2p3yCW1
FGSAz5QUpAIjpQf7dZM97hjo8DXPwKEXaEsfT5CyWquxtazW7TCEK78tLXrVOFSLE+uvtO9h8xmR
L5dG28c0S9FCTiewvRtKVyeYehqCrr8UsxzapU6yyvQC56FsdQv57/AB9LyelSLE24Fc5Gn1BuTF
QhGJ2doQvjEecJSR3igS9+dGa9+SECG1MlT/EhcaLWAWiePbgTq7k5Q2+sYwdi2zdqz22mK/vb9u
DCCk9xC/sg0f+vpvLyKgafBsfvQ154lDF1YCSCi2OFtSCazlQclmAJI9OmzM9xZvwrUbGGONCH1C
k6XJfl0DbRO++3mNRcJYTOeryu7+vFlbYurJJ5t25ebJHNUDsd4SgpHGaTWZuyHiHPElMyYN/0S8
t8wtK1ZrUIb1pyAomKEn8jd/ZVl56mCuTuSAggJC7wyHZqYreqGs3JA//4JKGm0e9rwLKvSgADna
n1I+zRwqRZAMgEzydVhKq3CGVMs6fxBxRKbCAV/2zxsXZ7/3PwTePMpA+lmDWjZkC0zamp2qOqLb
q/PPBPCrj4t+jOPRnXve7DmoVHmLzDxVWzYCWYhdPI+sFa9//x6YuAG0Bb7hRKNYSlEthvhhhc2C
hyoyJJ0dYNXlZtnm9GGVoPR69V/BFIiqK7fxnVrcWk4Qn9b6Ti23uTd1Rdz6wZL/8mg9gk+WFfyf
fVne4xrVeR+ME5ocEPXXiOwIPWOXQJtwHCqpFbWb5Rcge0x3bDQyETwFFDpq1iQbsj87FJyPu4BZ
HfZ6YUQbyiT1toZfzXqeC0NjtUEzVKN70AkT9ozv6Es3jwP0n1G3HyCd+j/nrf6KvGMVRBLbUdcj
2bJnTBThySQ4o2cMwcPGHKzRI6+dSTdYr22GpAjJbTktUGUIIKVASvfj2fQscP99WwWzwPrfX3f/
4XdeqYG362x1H7oWIf3WdoddfevteVd9hAjC4SuSLTdXxPUDw/BxqZYpl6JBZiOEZKN/dmC54sju
l3dKUEhiUIvghAO+lXNfmnx/6CvVe1pj0s6t5Y67r7ceNLLa3eMZo5D0zt5zuAFKskE+GpI07lES
UmWEbfHa35e0aSPKytRjyooe69GdJW0Ss5cSmsMQ/XrEUaL3qvNXPE9DPX4Yee/6xpzRJSedPgt8
HozzHi8GzSAZrfnRhkOjdLEj9G6X+7371L1p0mNSFvu2EqK/ukuiq7Woste1V0jBNn67ISgGiQsF
LyESlrypK/O9nlA/aV5JEJ0HnPlyyHTIYA0XjJSonLu5kRZE2gWbzF5IeN03ybwwVkbZh1wemaao
ppK47NwKcFLOM6+x+9aE/3XAlEwrzxpUGaX8qmde8jwsxoRrWTzd/ZHkEQ62PN3BWkm23qKjqBIR
9ZYsiKQc3hXjg1mnkmtAkHXS0rGJ1P2xLPHV/dmWBqFUjHDQXioFR9VwvzfBNnUoMBDNPOcIrsQp
7CW3Ps1rz+/FcJS6qFR99Y/i8s/LG/zDJ00kgk1X60vtrNlsd/FH7WY74tsfJcTYU6qZluxIroYF
7dbzEQKC7LZU3vrvvWMyfFfitOmGl2gVM0vU+pd6OthV3FsgSmVI9a1O23W+n0Kl+KOWUNIvjHWJ
VVZDqx6ff+QkbJrVqdCJ6obmg7LOAGFfbcKXuUWPyVk2eZY0bmsIpUW5cC1iQyDaWTNWDMzqx35z
ArJEQ+lKV4ZrWl8NHZPjMkCBEELQnWuIlVPfKuc9EM0Ie9QqmTh++Px50C4iOBRFpGn8xmR9ccGf
Y9hhPXUZ4Dzbtn2yc/Z/qiIowCW39jm7gTn0D2i/USoJVFob7YjhV2HsN+L1+RFxWzyX7iIlJhN1
Ci+NCAxWTWVd4Zr4ARpiFsdQKxXANVj4NspxueUgbW2bkccBGM+b+VXJTWHSeKJXUKtrEEhsvVOK
rbEBBJbqTh4Mndso//A+LsK1doqOwsVw/ywXRkIOACFYPqSn8+kpXGGucvziKSZBL5JdMAaS6r+c
pcIgEMIOtZkyStLl2anxBKoKFRl05e4x16mmgYMD2h4w9eCeS9jlvko3TbTqHWCl1iChiXMODQs3
F0s00IQThz+jaqeSrV8uyzXjlwAcsRTuGRFHSDn1MT/3WBZlxhPpd+proiW372M17bBvqCVE9E3k
vkymuvHcqyhsX93S5H0+/EVTAqjZop6HMNFq5Y16EQ2QcK27hx7IN9STHXhVEXJl3cChm2ChmxLE
SIgGh2dI/zL94nOa6ap7Of5yUYqi/eTVBopGnUXjuJko8Mj42whbGFydyhLleN2ILNrAmB+DCU9m
eIfngHgJi6DbVByqVr8Y+e0JAo7VtllOhoq+xGBiFVB3dvsM60QloPBQLj3iTSCujn68U0gYKlxW
AwpD8alV5bgMIISQlhvPEwF6tcunDOwRXAKxUWIIul+KtwSfXFQgcR4rZSlC0xa+aH/mKuFYNbUC
L0uO+M1FIihzNrjDyEz+7yi5GVDly6MUMa0Rsg4qNnpZ9eGRzdFs+CrYpMU8hfcaqzNn+9nf65EL
HHtA2spWHm2k+oKXqJiUKPWFZSuztPXhRIFerxpU2WgfCkTZbyAM03707FqeUa4PYJsieSKLl04w
fP4bOw2sUdLyRP/exhulwAiAal2w4oF5Wy3JTBm0j+I5D5aZDcutsXu8OtYk0769CZBSlGXRrvnF
2v4KQxLUo61PBHeWWjrMw13e9dyvS04ljvA2LMBI6m13DeXuiNRuzaSedowlfAveqIZ3paWaQFjO
8XIKvJppWR+qDa/xgi+rrS9VJpcF9ncz4fkjE/hknbV8+amuRaujFymYma+krEOMhPI7bkJKqSIE
GAieyY57yiyrQrRuyxM/lFzHv3WLeG94Plw2h//zUsE7xylU0twZllugbRqRwaTY9GlP747swvTa
C8ScY9XfR/eaD1TlszRiVdYip2yEnuKcpL/d5k4QY2u3UVQFuZzHGV1kCeo4pxF3hgRz8Au95+rn
rKclq3jRxNEt4x/zR3CBvs5T4CQvsI2HWVJOLS9vqYsVvXKH831boHhdC8/IpoNSWQzt1xC1++Ey
nzwvEaRch3e2WrkP1/Utc5owr4Hg2Dc/YE2Xg/iSSDZYEc4mnJNPzH5Y4uWnfMf6MubW11owKjb2
78CrjpYUtB9z5mRJVUWrhhRxuzOmWsfnvSFC48aJZPjq1iFI9XLL1hlezrDE2FrbtscfuyvcP/ho
FZ5pn8s2tJpjZgp7gHjRScI2gnp7iiRP2ZoZ86T5qh58ROJ8GkXaV5LSk3hW4uvqAYy1NjbIqK+T
VgEN1rs/r7G+RWj806BDkpKxZcIR/4JPZJzWNAwxo7pQXxeg2hjLg50ctiXsn0yhWksUhxGZURe0
YFCOVYRcwPJG36Wz0QWKbeajelzul4xi+llJP+EWWEYOE3wLHDPqHM8QW4Aq5eRmY9eWsWfqTH25
92v/HS0NkGMruF7AbQDTNcHFPaSQBrX4HMJCkj4LnHNVMJbPGf4a4++pllb/a6ovTOMIbBGDBybq
0MpEpKtCsT1Vi137mY6m7O7Om8IVqTlCXJ95NJ5Kk/lXXOeNWZwMJo3Wwk7t0B/T4ZX9I10T5zzu
N0UWR5ATqxmX1pMq0PV47KitqXvN6Czjhhbj98HLHRcdTgCtME2NPWhur8RWTtTSAkHOSxOtRggQ
fPjbFj833pRODO/76dOjm3NP/F5LABWBcKn9AmdzzbJvtheamPXvPXzJhcpR567hIUud3XHP+ywj
/sjHG42VjAg+Uf4+S7SIrLuD2akTbCXaPVUhnaXERJJzC/BIJnFDzn+wKPP8HL9udMSBbvaavszn
fBn95WTEtMAm6jKRWQDmT1UCu+hR3/a32Kpp3L0BJvBJ3C5ro36ZrX+tRVQDivEKY2USFvlN1l5p
R+pFCNQZLiu1PW0znd8Z6IAUxt0ha/0pLLSj+qw8sscI1LkBl3YuMcte8XwllTI1HzO/QQdrDQYb
wUt1IZ0nSspCxWa7pT3TPVjemB7gVwRh0uDbu74rXANGcUM4MUV8/5q1rc7GRereaiE8A15BjwYm
trn2ytOkRPwGl5DyyfS5/1SUw42xlRmK58D/WBN1GrDBSZVn2fDUf58Bl1nHq6dInbLK+/aUFu/D
BwNoGoZ+MGL05lOCaJS1YP2CcB2+eqBfcyTMqAQHyWlON/mpmEnVvNRyvKMJkIyiDip92cjcMXPd
06TonZFm3nQM7OaFtObW3c9HEVqtrB9vEVxJ/+ejNDTVGQKUsM+X5CD03dt0tBka7j+8uV1rD169
wl8gZxtiOFG8JQoazfkHO5PNHj8dxufzFQsXG2Ux4tNeSYAuSvktPCUqZzpw3MX8jKa64emny7mW
foWBFEGo2E5AfaSmW0aIxlXvJ7W/WNciAb5EkL33XXRB0uF/ZmMLdi148D8XgRlofpcH+e9NcTCA
qsecBt5xx8E59AuDVa7WpaZU8bvM1eOArbryJ/hrdGYAx9XeDGvc0ZVAxAgPzE0cTRdlx5eU+PIt
1Z30Z58PE6AUMR+RVwachoQy8+6awBiXqE1gsrP6+oz9Ma6owZkQD/h2nZIirdK+KBiQra36ydXh
n3ZulNiGYWovvvZ+SCHIOHy0dAWbRU5ealocEDVJ25oJqNMl7JVh95UkzxzOKnAaqsl9jo1SpbqN
Inw1mLUIshRMh7vGU2/EnJOFCCabPQ1znqFM4CCPfPc6mRx5RGSysPEXDv2AA6GFkuwDMT87RugJ
2EYzl2+uAJxK50fffVRKsOSjD4kJScT7dodflOmhH7jh0091Vv5SZrvZW+A011t2+5hR0/U9CwlV
ATVgna7ftGcLF+dXZFlNv1T/ZYdKWnRj5tVR9H0in66a2HulKp5V9PxnyXjusieMcRdp3h7jShjj
bIJk3tVfmkpq/Qx9o3QEKyZB0FM8sPFASs9JkjT1QQOlMfuTuYNpNlbQ89xddgDcDbsCdrPQptyf
X+g1JkbWIPhWxVOlIN6JkV6UbxE1pEQfTkYMKo/5A8GRoxLTL6tyHA4KfoXbj0T8Q8WcKjnDiBxN
4oXHZKainKJRqsYATbzPNtd76BPrz+7TiORSiR7BsQ5dKupNP6mkucVwpCTuWOBPx0+GL4ebeMxa
M+MluHdEs0wloGuB2vbqKkWo4zWhDUeUPBrJnCHhaCjTHDWn0hodrF/iOdWPIB9rnhcU2WxKn4j/
SbLWIpkE9eTuRO3aJEF8tXA4eU84vwoI0PD00diMBfA36Y6IdNopbdejSeOrNErOB6bBoyXyEgcx
5tz4/+4rrfIn/CEQzMLHFHBdiCIDgn4u2jzAJCmdW6uEYye18J/3giImRnVE1s29QD90xLnt3OWC
yOKOnChopUz2Uh/6immtxpe+qekRnLcP+UH0qGEsaADMzLWtFFzYuVRb4FRsY4/rRfW9FCB6ROM6
6uQ4ybwKtQcwOb+HH9Edy3AEnf1PrOvm/ii47lV5WYTwFGubRAmR4UzLgdnAo9/oTVzQ1CP340lw
9Ai3ZGU/WmWX559rqPaQznYKrxFhY7oWLAvfoEyDhIk2hiExQBLIWzaQJ4S67Eyia8vkbdzHqNoj
lm8YJqjg/A69PBDsGNvoqsiuSojxrJju4gNe3LTqRqFjrtqtvFFi4oafcvGlgnpGSwH7QBBYscHR
jcUNEP8SdU9EQdtKTtTB+vIyB83Ng8+mTiieJub2Y/XRNGfFjjmBvS4QAr6HL5TY3RIlf1/r7Mwo
Wzjgv39kvmqu7NrDxZdigvEkjtQlRXV5x0obqzj3iYMgJJH5vMjhGygwoyhAAJCfz8fGqxCj7MjA
pKVnHQDS1HrowxOUI/pTj290cShqAVzrHwTHVpe5h0rnsSCdO/z6lTua61sIqCxiFMg/slqd/r+u
NGv/s+gq2EzyN/OLRUMWPYU7CdWcYmlHx1hVZ2mG8Lv/AEMnMSl/FgE8r2mu9I8b8GJwy02Bhs14
j1Pl9upqDnj6cItQ0/lGh0R02fl/m7hOfTTSnTfNNHJJlH59NO94aL3RJ9VP2T7gvXsYyUxmza1M
uW2/gh8Claa9/uflXY+CvanShbozH67mK9s8sL9Pvr05AKCvCUzLbFwCqrT/8/bSy+dBfl6rN+sA
Xv7M5eUa3E8B8I9MIqorr0rxHe0jFaBnGQij7UUS/rxHPr6WxwTYBu1STukNI0XXQH0nVb/p7e91
tBpqXu2Ee5agwMqFhUhKIKqot+Vh1zObEjuFZC3FSb9FIpHYLq7KksLDqcWdYaZFl3XvxF9PtPsD
WbvBHzJ7ton1rrwEDrMOT2rKfNx1tozM4wPAeAqlyxw9nha0lhjaGeDZT/1xbiaHGEs9W+ngNpxq
IIZMYJiiSbfeLr+WO6hT9IMjqsVUC9tMwVPj1wlBCi/MyHktrtb6Qvl511Q+xFQpvxtTbdoHTAdQ
FMlrumKyMYUQwSaYP3PuXW6iz1WM7CeLI/05aGfYCrWXLWtzB7KlHddDosbE5dDrEYJLXMa+KwDT
H4Au/o7WR0zm4wAGz4MUrEhQfjx0+Lr/e/oOo2CqujPusA9aR/pZy+mgpBNQoCqM1Uxz881AyYcz
sYxHVZaWFVJrNyVqAmBLiRJmIquHYW8V7tcM7XJnpW/liOAG7U7XPzYDS/jKiCpV9oKzM1YTbdAs
7abtyRWv4v0OcHbYYZpEX/gveU9m8uCzImq3oyd4tQrnedymlAWciiYIE7Tx8vVayTwWIsYZPzRn
XEeFoEqEHHjiLdg+G47ehE4A8tjf0CZ9eXjcvyDeJxbOYcDKPrFIOIcw6FQNiikwiP1oZI8t/8Yq
NWUvOHzxCDrh/DXH/wsQLgPq/cJKmiAFdpBD5D5YGvlna2eCGRH61bNHRedX4lwPqYSLpGDuTqqN
ey336q/CEjUNSdqce65hkL1/ZDf/eAFdOFevUvFOFss+C6sDgx0D8Ye7MsUwJoQZ+kBBjc4+bjzH
Vs+HIrJxcJkJAz9UE2yqXoM1b3MTsaDQTBum5k5yz2QSm8FTdrTX6Cd4vxvApIa/qOUiFPZkCUns
9J8hgu1yJwa0W1VbpQXbUJqjd5ukEr3DxkHfdxpb6N1a0JB3u1TvINa91Ff8d8GOIy1viQjX90HH
OtoHEUm2g2f3ddtiBWRKp6suFD9CsP0caReCGrlX2m+H2GfgBzOW1gSxwYKsydgmMmxdhizQryF1
PKvT/Y2aHGt1+MQsp+AxewYeQTbzOs0pvSziBa7eAfB9jXamKaKURh5CiMzL0IV2N7Cv0CCtKfdk
2OXX6cIcrcqyju/0F9/T8OAdifUkOd84CriTFo8oo5Foeam2vezAzS6ov4d7Y9FdoG1X7sq9G125
T/sYFs/pAtQYLDmpRqHd2NDBAk+5e/HmWSA1Rqdet9IzQrWqsYd5arxgixs1cKo8I7BP/W5V5YxO
txSlYljgx+1K+B713CCgIiXFwctwwQcyyFKl3Ntik/RfKu8I8b3cl1NFWQsUuiOjJLUqLVOf11Zl
XvQOIGFyjYCoclYLcB7bge78GlLDh4jTNos9LK4BprtKeSNCKX40QEsXtqvK0FVK4OsFtdNWyX3f
dWfLiMRUKoOWJL2kTlO5q3Foh1P7uoo2Jn2a9mlbFT8l16xtS0pKOjLaxdfa24vJjUeUcSlDZTws
wzrJ4Aewz4cgKJ3EIVr5yNR6glDn3gmKxbVZYdu27ZSHCMK2Anvf/Y+qGKoU7we8Y83DnMeeV7wm
bRo/bJl6GBkuyadlkuLeZMAowG2/qlnEbXg6ix1igoixZeIYNqxjDVZEIOkTfQA0hPvXhtVRT7VO
nXb/wIGvhGnf+8f8a24Xcn4nYV+PMlsEhS7skru0bW7MYagV+vJvvI4gkXCMW6zGVl5h218rp/6B
BXj5a0DSUu+f4/AJgImOby5wsVMO3ltbIDYLnkNZvloMQF4gdoL79NrJCVHMlrVRtSnxSsHmf2d+
Hs6FxJ6PMxQeVZmif+5tQKjKHgiWftANkAv6yJEeuSFP/V8/Or+hSGONoWuLs067SFUcWvFG+7On
ta/708nxWL3ChSzgkC2VeBWj8H5Bsac8DnKDtlVEr4d6mB80Up3Vr9PQGiy4nG0G+HvhM9byEhsQ
CRWx8BiIR/wgcZWuckmXyUZc+gqy6jBO5anV9daYw5p78qU0BBoJPk9oz+TXjboj38TIZ9kOFBjA
Ji+27ALsT9maJDn6yR5vz3PVpd3UHcfb2StezaduE9RWe7/+77FnLAVFdJSh55fP+3P8QOIfVNMk
P8ZI3IQz+b2mBmkDrVojnEv7nazUCZIVOBUkGO5xXwR6P1Z3saxXFq53o/vpM5z4TIvNMaakWlba
faOfKskYmqOcCXE5Dsr+qIkKCyRwjYg79Rlvw1kNYpOmylh1TxQZCoorMeuXUBBPzIpy0VWbbeuk
2OdFRFh3MuZq0rgFzmtLNOMHffLaxyJ52fVqBg++RiF3BdRMNDYzBanZK96oQakLPXNavrXrZWB0
yX55/YIInzv6ZGCas1taH1ZghhOrmsjQwlhhXlTeKq9f8sAVl8cWU8pbcT12HoqDlQTVI9c+Aci9
u9QxZZ8gzFnkxWXJ1KS+bSamveHqLI72MnKD3vryMCR8EEs1mTwERiIDfQH/jEu6SDkKbUr3iwjG
NUT52AwCOZCmYuBvxNLr97QxWBiLO3DzY93eAFuu4DomE3ysj49uj+w5U0J6xiHTP7biv6uqUw23
YQw/4UNYnAOfA2l/BNg0eq0IbXQnfIxt7LTuNpX+fZAgA6ZJTHsqkx4zUIrFD41GAhaLWFVoq+x1
luHfBSZA3JZOVwYIzVpYPmsHDc1r0KsqUqAeaQQA9c9UkgSW37vuy07y6NUePQTh8ELO2Ewooc7O
EagYG3g5Ks5EXwmoREwv2EPLO0Nvl9yirvh3a2n2+xGaCPlp5XaxQscLFhGowMeUXecBS0sT8UZn
zsiWbgSEj7yfH5fJfvJH1NR5fhxbdErmNrP1BpFwpdlniDZoe8yMFi39TzsgzHtkRHPfAvkEBCJr
N4bS0DuJE7LRf1sfxcd6aJ0fpzhSe0dE4PFV2YT/+7GC2Zof9q+ODMAghyzLAwaU8op7JrLaM5LJ
34q9xbAhKY0GMqHxO0g4LvicGMh8S7WTNr7gv2uRoU/RYV2kx2HqZLvd6v1bJOTjUOuIvzRYD9Qn
0JDwvotKLEORlNV3podNeVCjVVXlXN0wEeRucSaM5Ye1kYZnSZpWN+Bp5iGVY62PhzzST9ayQrWN
VUWy+2gJW6XM+3RocYAe1IvD3V1/uNCF5agdr+tDRdXl75U0A5sFcnTdgIoQh8jXPq6G92/h2Vm3
fuEXeQdLDv5O3O31PDIUCLSpHCvuThfsBUjMfgB578NPFRKNsiKCp7P+b6eXHK9h6ljmoO8G5ix9
OPXiwr/Vk7MF3nCrIYvrIkXJGVuRzr6UidOPLIEX7rc7e28MqWEIJrMNpyVCyUpEFJnmLKxFo0YX
SE8sTwODje1g1dqfTX8AODu/Cum4NwLT2agqzlO8OQco5QtdRvAvxSwKCwZd7cuDkNeScnkFKPuE
ocV9ykOmDNjdRXVNq0lPW6JHMn6t/oWZPCUib2A2S21fmdnYHgRBofPF5dU83rhfA9ADiKZ5raEn
tVM49QXYM4ykBFBOmjae05N4PX8mjzqLClgMzthHy3UYzNPWXFAQostrdgh3BUnRNmV4XH/TbF9o
Uexvd7MYzwOX7rk5bVtlZpKv+pPw6UekCd3gwlHSbrJb9XK9UFEaItaq5VQ8bI9+pMKcJlEqUXjT
3hHK9CsoRudn69FNOwuwHZTTl1j6l8HeslS7Avmc9jz0Rv6V6l7K7nYBpi68A0s4b+ikENnhnUz1
ks+q7FJShJoNQd5MwhlcDape2kY3Ie3rrfROv5X2kaWHGsxo5sxjyq+PQT2hH1MtfdRyg0wHeqxa
qq0PHhSN79bLnwZiT7GNRN2L6QbpLwkGsqsHq5HPfU//4z0PXGCAAoEVji7jhYrBpmHA0UqofvmB
aEdZFD/NE9RQPjHhNvrWqcCSl3w7t6LnXKIeHpgmKNMkbY+6vAC2hT2Pwtyk3eKXCK2YD0VrppG3
1XU/JuaAhCAQ/FNx5ujIP2HZWKXikFiszYbBGffYQJcjuNyOAlxCf4ANYJc/85E4hl7wvQZ0FYGF
X8RjdscnKg/IF2+8EOcnVUyuKZFc6RfVFNX8zywB8iJ8NpeovcpB0LG3b1KVyYfYhvf680xKGw0m
e8rfhdqoTJjC6006PawMfQq7GnToLzK6vuCsMn3OtaoYL/wbz03d5Q3IsLOFJRLnrhuIXugB9NEW
KeFIi/Nv5H9F/XwOugkV/RxtK/SVC2nR0Bl4PDdi1Yef7rzR7GVdwj9LjbxG3rQt+i22BeL935Eq
Yj2krK5qTThomUiYjDzGczrj8Qx15pj2JHp4HyGa9Lhb/0/YxPXlbEeivrg3D33XqToSNiwtQECi
wDyHFc4jMV2AQsMbVB1IsV3CS5e9dXCcLLMmmZX16WzwEqBPBvvIqvHuRyJJCNrMp+R6ME5XlMZS
GbjZthjPyvS/T2WDui8VLEWbvU0wypWPX15YygdgUnF8nL7FG7Wyqa6s0T6/Rapbz6TUoDUXZ9nH
B4PrSkZXWXyJGUp6WiX8ABk4CXwXQ7YPUUcd/f3/UOVqgB0GSpeyFaVKXQYFYXHndcPdMgXtGU8f
1+DTWhuN9io/n27SHVvCk/afYP7URmjTts+qkRbeiBqV2Q1NpbbKw9pIJBLshc8HYi4xdWymioMg
TuTgU0WNXEgYILL9/P4jg100CltC9wcuAroBqI1kBE2ZlR2iQLLi+06CDpehNmPq7nHfY5BlyRG2
YWv/xO0ADX6/lIA196sce6vFEROX6UiXtOxvPpcrfpTvhjErJSgPoct7p40KEERAkTQOrf9wmG75
GTQbos6BFRwGCOWZ8EJRfMrntIazj6xAmkmzTb/gDZSHkyLyoIiikrnBpjcuyM1e5fsNtptRkRzy
V0p+hAsgCKZFoIO6xtQRlcc5tXQHbXJbJsorDmAtB+1ipNr28y1j64Escyylrb5sh8K+knxaNY7I
NkPIiGi6Vo8YKo/j3b4f+80Yrh9DWMg1Ga953L82mWvSiBY/pwRqFiLtfHAa+lO/dkyuo6/xSZjT
V+AJstHLvrLx0GQIzedhzxTSphUPMpM7GJXKDvvJBN/tId/GuZqHpXp50BRsnQMlpMTkIYmyTQlQ
WtYeN0/BV9fg1kJ7zcdEIj+jYbGXUYpBCJTQhx50YoP0MJht6hOtynyk1B9wxQj55PqEBo3leXn0
Q2YAfAW9IZ2AvAeTi9RR8wL97keeeFT59lcU6Myu4eQmT5gW8h7y8mHaWC0Vhde5/Tnr52p9sBu8
i5lUNjBrTldMWOH2Sv+5ov4J2/cMRdOvlpoJYZgDdZp4xiSFMpeci3ReaDQFNYiySf3vaZNyW/72
RSO7zPOGTZjkaDV3KM0FeGzL/JZpnySyXPNiiOTMLwz5QKIg4JFBnXCRfv4rgyy7ucmTn/aDsHdg
dlBKV0spTehJ633eskEmxB1ITQ5h+e2fUKKMO2/tM2+ANe8bxrv6eqQOvMvppAXtaMow6L5TYUfx
PaohuLLPbZQdVZmZnsYOhXyPbu3DUz8g2ql/uirt0v/en+w6QWpPN4GP2035BHxYe1GS6YI4xDOu
cNVdVXaJxW+jN7paLK49tMPyzagAMpIeVhG4s9B5aoKGJPIEEkDxsP+/TbEZP4afeHQGipzfT80J
mWGsC9x4r/yVYFeO4lyJGKf10irzNqfIbTg/3tiQfbosV+sH5cOW/6t29IqZGRRPKYxAx4QzwYvU
MnuEM0PjMaTCKTPzhW7NCqf+dIXPxgqx3gxWu+mWWmDCuR8fucHIfahvzwMfqP6YM4BQFOQUIFNN
nv1n361gquF42kEDprlchrDQuCzM97gAHFgANhSlLR/4qCbtqLEGHC1wrw+gecR1pZuVoAwX1f2w
vo4SH0LHip8/BYHufY67WkPHa00zKeLkwXBPnXS08vAFp21f5OImSa/Q6pzFNI5eGEsslSehrNdO
VXcvVj19i3fgukEH3D/P+ClnD+E081hHh6PvU5R0ZVsQxJTiSXnAUL937euQewd2Vb/jgRCU8x/V
06gFKE9rgAECJWLLZZUeUYgp2GMi0KvcXBjBOiNspJMwFLsLZB4eR24CrceMZA88nTAp3LGJYzB1
4bLQDNLphLaob6EqsBDcl8xm3rEwRZiZDZUUP59MkNEIeaLa/tiX2tt45acvhPyJ9X5HzsZXcURu
DW/LgLbK90+TjFmJTLvKXtF2l9Urkw7dTgTqgSvxUIph50ERga9ysZdWa52rQHSuOzzOT9Bd6Riz
V8MWZthsO9yT/BVeG2OHPBjLg8HYafPwXfk+iSkvSpD3wG/3FvF0TtluXh63d8Viw1w3BXvQX7on
2CtS5FWz3wUh17GmvyFWmWgdi9U2ZOaZ0zcsSEQVh4DLUEkqb/yg/7bq14V9fFX47vW2RyATGRHn
vBSScUvyWfK2N+cHjfHBuq7MOP4gOweiQfERgGXNHb+Zf9ImQdDBzO4xqylWM8D95Jyn7vjSMvZR
GXNnJ7bePuXnOy7Q2nuruhQKzOvaSpXUyLQlyLtNbj02LZK1V/P8iTtglfKBWcu8/hc2FBBkgO6i
IKmcQ803cqNjB5AI8M77Eud9Y9LjFmT+49b+Tba5AxWBKBAsIizGO4quL4YkEQgjL5sH89s7YoQ+
A82FaLy7eQCBO3WXrdOhbyvo5H4/3f8lzFR6aekoADDdKKodSUQRdhCl+UcmfFuPGvVupGCnKuCg
BR3k5BfknFG/h50YjXCIUCOgu+srTtuaQ8IDZ5t0ED3tFlr+YLK/Tz7a9D4MsMe3QY390Kh2Wnhc
bwfzXR53FrHA5JYxqxzv9CAgwKmf0ms2ip2m8n9A7UYD4GpgnneVB1AuZb679DiUfxlsdO3ZtOYx
EWSBThQRmBxjykYfb2zTVi8dAvQnOea9Q0MGi3m1+xMOyrwSb0rXQOFQnDSgo3fC6x0LcgYx+Qcy
dciqG4YdPIC74rLA/Nvptll7YqZBFC2DZ8zg9f3MYnk9JRsEVeoa1ZUHlnCYnKpyHPOwAJg7jV2M
5BY0xS9YINnpDHCA5cypaKSrA03F74dUji7WHBYuD2T25mDu04QnNG5MAX7TQanL2r6j++GxyDxE
z7hljfdElnQzUZ65xkcTH6S2WfQcI6Di4mayb0HribYbi05BVFL69Ps8vHEftKCmoptLEJQYpRxx
wm4Eb3okjFtVtTbRtGqBhsYUzal+gfaLBzHGG5qMdaBM8Qsvne5jml4Dwty4NjnrzNttIN02QVtW
LZbQPTiZM8CXIsL97TLRo4miT0+bqbsv5G38DBTAAKWDoz2qFd8oxL3Ft97U5mnFLYYuMZgm8A3T
qY4TcdRfKvRLDTY2v3sYQOIng5Bih0MFHbdQ4cofapRgeIDvBqS0qjq+XL4PZRLELwW0ulWUEfsG
Mb0f0TPleUoBkCQFTqP6qn9Qk0TbEFCmY+fTjC6nqYzJG4mD1OJw7Ffe7IrscOHZsWS+b8S22Tek
jQfm8VjphQeAAQwPhOKkBM1IDPWqP6cfszzm2M3gvehfWDbNoCzimmdFt+OUWGRwzWXv6WHSHbxm
kkNOdR0DjqOtDPj/zhu3BrIUShOHBJ9OTni0480wwz5iQWPEDBDZdVtBmQV0YSoLGBcXAPzSQvtD
FIxR2IyvW3SInIn8wdlhtvdPkC1f2Uhb661dxyWJI6LxR1UbEkM1qfwbpx7VqkJtB3R/OG4oDqi/
4dmgU9jot9c1qdrsb3NHqRNwdYEy883X7jP2RDSXfX6PkPU2EtCgLMijBJk27zRWcyKs4rxk9Paq
aqhsAi3E0Mmxv2QBWGU0QVGvxnh39+/9Wp76VU9T460srB1As1XhimeuPsHcJmi4sFvEN4XrIM2U
mG/FRjGdqeabuzaFdgXk8z8AJ/nnLP8YzRHXT9jYq/wFGhpKgRBCAE3f8oCdz8dEzZqalJzt6kuQ
px8kSaVOiHbNzJQ2ra/Nh3NhRSUWVr9mVCgBUZpJ5JmQ2fky92t4xmrRukf/BMdL62TSwSx+4DIq
tuAH8L31uhsAcu+bbld706Ldxvpwm2RHBHppLam6NuMaxevIl560mqSk+8aXQqblofFgmFQnBVqX
URLHdhDvVTPCj4UBYXBxFzV9oVdvn9OK2E0IJEaVhTiGCZPWZfFZTHekfk9nbkeafnGEvdzs54Hj
gJPfGkwFvNRqFT2e5gcuF+Sw72+onLBPb3x5cmKTZoVZYVizWmTcroMc4ZTKvsZcwGigvwz6beYO
JzCRiJXKc4ipK/ZMmgrxZLn+QBF97SShZ8CFmfiEpZPznyjHSCwaGuHTykb2llNixRaZUaVIu1t9
ZXeM69VUSTmoGGJlEA/7WforyJgUW7XLM+XB4ZVLqzBXSXhB1mWdN0cuhyQb+/xOQT83BsnrnOJZ
XlkvHCr6Fv7p003vCfBW8+OMlEK/9bWoXGKNn1wMJucB9u/CqyzqWRH+qz9/GoX5NDvycwexhcG4
1j3p4jxtR8VGWAE7FfcxSRdy6WUb3FqQyJG08nkMQf1aq1O4JLElVrbmu0kNNn5sWsEQaZbQhh+d
xRvjd0HpKIoGzRl5u3qK4tXa1lzXzAOhU67oAMgTxd4d/Y5IZ1Uc+5BXN5ay/f8uSCUUvmYzpBfD
GHmD6sO15gH5CPwcHIGg3yvJ6op3OfO45X1X/zI1UyjEbqh/ZsDp+Sv9RZVNiHKhZTbvrEQ+BdXf
X8gk5oeRLc/UvU19JKMWddVNCZg+u415KggVXd1/mEKY/4JlUf8WvDKVDn4zE9Xf51SUqLq+fVB0
C1a6D+/5IrbcaxpsaVRHhhYxWzyFfXJYIlMC2vGHVPipI8fTNg7CiNba4D/Zc3EtSTOXNljDdQYl
w21bWB9N7yrV5BuSeyUaWy1aKl0D1pGlJvoO2SZWt4QLSUUfi/qMhvwwdA+FCAFvgMmsmTZ/ie+a
LPBH5fUd+StdPdzKxRSTGYUE5/dE5WDgVQQq7oeZb9o+7u6AThNzxEp/80KqvgEg4Jkzbdwy3gbT
3GsnvHYD1LqhtkNg4kMD/Ys67imX+VEYziSN3y+AIcfQHKgRHeSIAMJet7DMB0ohqRbAI6Xu2yMr
jMXJkFYfd4sbvqVg6gZXR1K/N739vqgpekW4bHdgZ6rqrvctxI6jhHfdRjm+4sJ6tx+y6YdMVEoB
5yRHywZHaC4it9MHwCJbrnjgOQUn0pgKbHSxbTbC0W8em1LOcSqGrqwpHPsfkCEnDyoFYGRfzpPu
SZioW3Wcr/pzoaSobf7cfAo1ok0w/7Hf/96nUXlCutaHpaiZbWGKRg6l4azq3twYN8XVyJUOQnw3
NqLjAOy3iNBdGjHR5Q9pXT+XoCWinRLq2TqpZXI3t264Wx6ZYhOkf6tnfBKmOQk9yTIdCPvCT047
EsHXEcjE9z3JQ5Ls4k90UYJv5k89BB66ox02PuQjQ4dNttzMB5SPPvt1Td/W8NGtyy+Q1h1mjdob
ncvvyUJnc+HGjBlUTuo7n+b7DtlWmwYRg3gRCq65HGyNQhK5/8MqzgC6mIHTn0lcGmCEyDiMXxF5
0MmzK2zJZkkcgqa+y3BJJbmdX5d6EHeIT2/W4r/WYHhT7rB3tDWaPeXyMWdUhGFCcCgkGPl+aVXB
HNnpv38f1fgkvYdO0/pQFp0CxzlHKnAW1xHnIRpvU6Oo1gFUJvENpAckg2CrUgjLl6w1w0rTkVcE
Qy0zTLUUeb3WGnS1w9FaIiPIwMvbIJcFL00N3fQymeRFKeeFAK37xjd4Dc4J06KbKpbnXqKKR/tn
StUPAQjbO0cfPXxQV9Z/DXX0DRHE2yeWVLUXWZj8W5uujqmLy3ab1hu612rV8rfd8+3zTeh3w33N
f6o5aAjGNfyOm7/tTwPQAbMOp8jXfOBHRbiJYpaRsg676+hOPrZZND3Z4XeNJjq5HmfXemV2nPcs
zZuSef+qiRVqntU3Pxf+mGvELrTbAl6hq4G9NEarY9zSlu4PxE4pircev1tzjuZO+PIvW2JhClUT
UZyCb5Nbkh59+qEPPIl5kePvfx0GxJ73EGGOEiaT6PmC3BtFTIAXlog60CE4s29AfJpZELeuWcyc
Fcq9Y800Xi3rybjSuO80aNuH0p2UnqlpteqzCKsbH/Bphagc6OIKZUGPOq/jM0p7oq+jx3F5P/Tq
jjeGZZ/7dKj59B12Re0h4lfLo8e539x71ju8sSd3YYdrXMJgIR6XVKnXrap3kCAbCLc0Bqi0DUxw
8XglVZ5NV2sudDTgsSSaIL9NqKs5pboijy5LkjdlhtZWNuiWwcGcvvP2zr6pYo+2P4eHuwPG6/2g
pp9i6MFmf6ETAiwvhBdQrnKbukhxe91OGsTSLaNMAAHYa9fFgcw9Rhfv3ra3XZPv3AxcgJ/X4dhB
MRj37I1eMGPrsK5AJ6QWns5A4pn3FSv09/ZPEce9hgfIOlk9+BiaWFpbbxlsZCDC/XaDiXiB3AVN
2CAovu94x/J/lXGTpIDHTXKrXWvhkNcPwSsnhMIvarf8+eJ9isZXDqYgywrA+dHGvykx79zbWyCC
QdYm4x+Sbmtwe/GXdXSX4mNIp1NPM6+6wrfdNF8i3/aGMzGMX5B1wpCEGpdTsRcpMZem8eepczND
CtN5mZ/sWPrPuHvv9+nHbSRPbVnmxEK1pQA6jL9fVlk+c2wYqV/SSf2FdWzqI+LuzkwlrnMz+Ywo
V+2a0VVMXIisD+O/+kaEVkH8c/+YAgtnXksjyJD3z97mLjQezUnrN+iEwSzxwsuR8+mx0i5NTbtp
8FjPJO3B45vKPSSJiN/ZYcaSSWxkHivWjBtOSDv6mzEM+98cpgxve58L4Cfc8RDLA3hRDfNxXUvC
v1qyi8Iew031SHlwEQa3QLHgMITpYAjyI1zzr/0tSi8EBYqO/gNofoE1rUWjZ6Zj2jF/yC+6+99S
q/LNe4J7IxeiYbjMVlbZpaL3I6aPgZiEIeAHcjSCWev0mV2+ipfB7TmB9MgSE1zmHXdiDba/bGYM
Jf5RTv6XWJ+pLE8xrDTMP2qjq7Yu9gfyVKamdRtiXy84n7ZMY63EhKOMCedPDqw6r7xmgkGtdHfT
hGHLO2OHHzYt3ZwYQUp65XBrUdka0dGndKgWSylTCW8fr5xCOEE2aOCoFDXTShKEwyMLoplWSJr+
PBHwdQZGIw3wF7ZU0fol+LHQEwYzFQZYT9Poem095FFofjkvY0DC3hLjcXWNXDaWyqzCUMcCRq//
5Bl80FP3MYVHrkXOgIV85D0s8eEu+pRMJcmah0YcmSP/kxOKamU8L2rORTfmHzoa4M/q+ilOvYLd
Gj0+Sk4fVxt80JaDXJVF1suO+hm7Tgeu4sSDbVMGEdEv9E1XbXR83KXWtiur7iab1CQTwtiHNI+Y
0QU/oR2Gf98BGQiAHgcmPWMhnpRLQLsvPZjDjjSpPJwXigUMfdcDWfITJ0lLWdjqk2aTnkgQtjdS
C5B2TdILn1XW9U3RoGAIGHTfeZ/0g5HtyeZ6bjFE9mJakqs82SkX7BOYhuJYv2qrZewGCv3wqW+Z
pBEsqsyT51j2ot4jyjMQ+Lk+uU7w5Y1VNsedww6QcXx9EspkaFi32hjP22wwx3lPdGLzDHWSXcjn
3YJmp7rI4TTPGdqm8KzZqF+kaO9Bt8gqcarW8KkhVqQAC2r3NlXM24ra0MYTDsoStuymmHBpDCOa
w+uqJzCYtYVvOLKSZFa6FGXaFs7CMUlJ4rNSjRP7tAN8ts7EWcPtRXSSSIKdPEqjzeObz5V/O6zd
ZJlXDtedpuH+yON5BHnj5HE/fXo7S29DOSc7KfE6OuZJ78qNDaB/TptaE9sn1+eHq/rPfLKMJJPk
/ss04zTIutcN9Tl+P/ugvUY4R0hj0PxwwcTbxypGcMxgFRUS0LsaG1BbizBNqH2heZmFZb2EeEB0
xHaQ1V5lqSWVrp/tJmPWuuw7BI+/v/ENvsZqr+RLPVDaKN8dnVNVI1Lja0stWs2IslK9gq78h8CR
rMn0pDsXdN5j6RVBzyKo1AcKYHqAksaHV3uSrW33h5l64uJj97wL5zZl/Qr6Go43C0wiM01d3QRn
4FJLxP+lUSFbrUVqqAvbyGuztYEuW4aLqFm6LQIuEbmNZQQsNSrmLdwsaf8sQiaramZe4sg5JU66
8R9LT8HLTz/d1pR+4Cqdz3S9/WpY0UazqY50CtCnLpBz99QkshFKkTG87x6V5cQVkfmcQscfVCj8
DoOkiWsVnLY6PsF+5nN7CITculX21/fDa/JgcQl+MzK2HVNJP3mEZFsp4zV1HJMbsomnA+n6bWA9
Z3Rtfex3ipaGf9TdVGsCG0nVU5gBRfceZGKi6szRcY/Tlu0tiitJ64doq51r1usFZiyzilHZdq+f
f+NUndYApGqHdNkG6qFBPWLE7qiiBuYkbMgGVTNGKoqNr/Wx/qcXehIZwfSqIIcqpe79JHnl8om/
f/lmFxKuVJUmvcPTrZeMO6etvE9V3axnLCzlPcTh36A0VqydWVnVXQ4SpDWopXfrDubYGGy5E1+3
8Y0XooBXBRelQ4ighXRURRycPVPQFUCLbxFXuQq7y1O/W/bTPDGPWmfsuGk9lQC9O8jUDIavdsZO
mIbdbbCisyJRdyl3mMiXlXum8blY7FutZWXX884rys18kdo9aXe/cQG8rxz6ExrWwCZPupsrmkGE
kqP0i8Uq2eQcoZXa7A+Bt+UFwwhGuHepTyNaOVkr+oD8/k4D6tihFDYbINDG/wFF/q7KL5OljGDb
JtCiNisl6YUkxlq/QMQD8FydHXdK3xvq7tizMk8nf1UBs20rKTZ2dstq6A3Ev0F77LkcXy95KHqr
G51aI2E6DJuRL8nU9RjTqzOrBZnOCI0d811d7Uuwg9bPBrW9t/IaRXCeGRn7EIgd5fKyGR/gd+b4
2wgn1Y7KoNzxSBzWdR+p71RmRfTrYW+gmvNPOUx0Y750FFfaUePZger0QQ8+JaWBPR6EvH9RG2xZ
g8buh/hfehoe7sFu+UsdDF/hg9CWRDZtfQ1bjMLbJhm0LBeddqQ8K0Okz7ggpd/GShn7LwT4kpk5
HW6oMz8xSijlE6zxGQx7HgH8RHQP/aLeVk1gqx8+tON5UX4dR76B9HhdwmkQcN7jauJ2Wac/W3Z9
YFypAbctkbzQfJmqA+IA9BF9G1i7Cfzs5bWCpt7T23E6RpRcnjNQoYSkTPjcn5cXFO4lWksPhq7V
XF+jyvF5t690pmSMC7gxfnfPS62v7MK+zPcPmQEU64YxShyXxiEwfrI+Tdt3ek8a9nGqFfw0aKMb
4EXorSjYG5wVrGK5EMmDJ83IC6m9QeEjQc6AZ2HEPnApIJhsHbMbO4CQo8q8Sw+WaW3gmS85RqZJ
RyLQk4kjJDxJ95Jt+vMJ6OYTkvHwbheL7JK7LTgN6gDqu8ueKfnafMR4aarbu6kK23xSAqkMQTom
oWJBdWP/7gxpQI1sgO/yn+ehKTCpJyrmM6elTbsNeLKuVdmTOeCprBCgawUnzU1G22eSRlh+521T
uZ7r58aCm9zcReIbsGR+yCIgl26jgBTXtwaPMmtjB6fpniHeh/MpbbqWffRw3A2/c65MY3qSDam5
jetlgLGFjvOIOXDl7GraJnUb43+OMdUhxzD0pqL1cwMe1KKdBINGFc/jeJhTBVTff3ANmSymcp/e
1Meq6Pe/hoN3zNnEt7GpNrXOfUWhpCKy6JE7Vhvm5Vt8bp9Jzvai411MKQ/OFNztGdtVb5qqzFIY
7FXUmtJEm9G63Dz3qcoDjWltGqCbJm1JMlRo4Xvya0HLN31GQqjWZGdteRJvj5RuvIVXRO+TeCY1
JKmOwvoTxh3yQ5A8hdnNLJ9oa2qNQ/WYxfl+ptD+NClA3X5OsPUvlLGaUS3bLRj3rDdtFaaRms9h
97hOLLAHGo7mE1UGed2DltLzG2O7U+REICs+PrTpoulYTDUu1k2SiZQ4JMUeTfiVjCdwQ9Eogmuf
JJJcB6lv74Sriq2B2lXOjJhDocHgjFno0ya6odubmWjzPmCDlt3XkMw2CDj02pnRtXZWsdWjN5AR
MS9Sr8KQRNVbE5SOqDA2lsXEOkOiUZaaf9EmpkU/yQzUbk0BOUYnMeDg4AVP1XQaLLRRKuCkfyLK
cQSo6GH7QKN7dm2aZwAvLcUY9y+CCe8suOPWiRRt0DOSg7uEFPAVKkkVr0qnRdvb69Qw1nWxne7U
T91KjYSlXLpgMoKFfmVUDVfbjIVd4j28HoMUH03l+34TZ4/TcNqOfoxF9xvURRabubY54zEhvOW5
rhZtPpsHo7CbbWmnrjhehJl+eATZc3wO/v7ffbNSoqOz+nHheTrd0lST6Qo4hlYL7vkJgL63nLS5
1/qL4GGzfE+8DDOR9giTF8c9LSd2lbpTUu/lsc4SFuIfvkDFKxT6hk1SOdVUbWtpQW1MTLwDRidw
uGFWChsVTrAA2LieCfLj0aIJj1e39gPbzVjO7HEC5rWh1rzgnuhtTurlvWkt2dnNWE0ZgJlsGxLV
C9Tz1N77ZzSYvDu/7a8jbiYCDV6uPTjh45DOdgzpnzWoUOzH38xC3Ndj8l3csgVFyXlIGNfV1RO2
c6wLW964C2EzjDCX21L8+xEL3tHgvUCdIB9crP3XRR6yIYBWP5CTwNUbXvLP1/Y/CcQeoWr2vMVo
OI6JwvzwOUnR7RA4HJggNqe25mWNxulUngv8IJCEC7p/9VOh8gCcHTIJ4yEIzqlaqrO6eSHNxfUj
WF8F6gv0uXzMazqBw4gnJ/Jwl1zvqr8BYh+JJe7IYh49Qn0uo8uG8AGWJpUQryCBBV1gxmtwsGEn
MKEMTeAQvxwIN30074mYia8aGjO8AapsDhwVLH3IMktSppQvuaSlaE19IMXbLsPgIswk8JabjN4n
t9LRlL7BeyQkwI3uvnTYppu2r30KNnG1VYACWWrQtGTxhoEXiltNX4mJOlDkqz/2jm0eGN4AaOvj
7JPxhRkdqDMg0xvXhY+/hRp/IXfYwq/KPem5FHeuJYbck2OY45M5npnmMgzeoCWzVrfa0xVZs3Kz
2GvaWTyYNAhG4atJ9hmwzn/bhZZKC+g9nDY/DL3b0WGlrNytHa7vndsiqBrbAcIaBotnPMiKw1Ik
A+NWGPJLnkdm+lOd74JABw/rnICPLmTqzeD65QHK5qtnIF/gOyapjduHRpH+Fn1qIvDWysWcho7e
DNOuetA6iXu7cNNkbuZJlvSkm/03qHPwfn2rXmuVpTiGR5hIInB0NmCWm1u57MJr4OnDQUjOtgH8
KnJvbVwhTgJg+L2f0E99Ni9kt3zXplZBPqPwVtnETw4KmPwAY7JZ4xm1S70jgjZPKUP340VeFJPL
jBj0X6ziV6X6bU6HLTwFY873n8gtKdzv+mIg8IrF/NgUk9i+gCYdTpavdszn2YtrM0/TSYHbHvv2
qOtttoo4OZKrh/fezmXoFyFqByqij83owW9u+zUt/o8QZfQy7f21Max5a98tBAUko6fg8XFtJsJ8
n7QONDeb0pnQBXaLbfPj0TbWWqfhEWL37bPvI5SbsXfhUA8dt57MQuSkSRd9NjJfNRyhV/T6MTAs
hx95W8SEmjdhraqyj6zUU+5c04I5dD9xcb2fmEGkCgfKet0ybhqYJpkMTqcr9XZrUd/i9sOGlOTK
DBDNLBv37K3bDw+uFIHahcJUiq4R4wnFrjDZYtlRruF4+NDhci2nlCWedYxF0yJyBPi062PmpxXb
P8a7d3wSIeFxRt76E2fMEsyClBBvt6X4oXi1T/IRmAxhjiO+BAVJwM52K1N89t1lLfff+MxxP9Ur
rfwfIl+auv8vjmXTpRsma6gEJeU+JakE35/o47a/LS68N5k1fp1GMRLkudmUO33+5fdHCsvrQnm8
F2/lW75Um7kkzU9+NLfALWx9rf5iA3Jj2qMcH9BOWe8tKr5wetWxcHCzrJvms+0rLdxnBmxXNGtr
mPuNZakHwUZjZULy+ery1jqP1UXdnrgc59FHCC09gbBmtKZY/d5vir4I2e71mv1WeQDfpcJiUEVH
ymyifFdfpe5dFk0cgXGh9aWPU4dsYws88qkrLZo0+bMwskzViLz1o4nj7urvWHg10qI4FppqSTbN
H8yW9yeoX2CoRN0rrKdu74pXWRYSV1/LOLh9E23egGTdiVdDTavc+efk45lJ9qdrmXY8/4H3TIna
p0oO37D1K5YnKKtRUwVl4P+IryhZ+z+UUkYgSpNy0Mk9UpnhS2hLZ0YLS8wp/E8lBk/cfAEf4AV3
tLLEYLskiTLy9oNhjW9eU9gJca4DcJVGrtMPIIZmg7QSpa/jgxRQ1ermx99iqKAOp2dC0fSXKsbZ
79j14uuvy8/TDd7225Ug6qm/0mWEsTZev6BL536RkUM2tu/TOI7tTNhPMZwCaEeL10YV68qqJcqZ
tjdy3hGJAVWYeJKmf7xG3VDizZ5lz5QJJaMxiG1N54CgiPGoVPr+XDvBNs4owYGtqMrbh62XZO+u
1b+mqPIlBjjHKVuUwii5wzpmgLuq5UBCH2SBGMOafA25ohqSTmL2Svz80yS+wVL0bIVswe/gjruq
oqWPAKge44t2EjKcuMD9/7zJ1e7Cne2afaZf8vM3KQ2gw3I1/cKvloNpSHkINhQ8tFPm1IvPjj9R
IrnozaCRhF+tAYQ9Vjy87imlwZKkDvSEsqLct2q/dmWTHjZIjwvut/ajfQXme7Ach1unqYldjdn/
8DzGToMCzsgSP9P59zUErGo8H9asFwYmtnlmX4pasJJnw8+VQA6DrSj3ZORNEkCdSjFBxxuIN1i6
qRKUoF0oinBv73KlvW6wNn4uH3CRl8rUpPqRBo2o64e0tS/NqSADQ4/00Vmr0TPJiZ3ETcMsMY7P
KglS3tzbnIpUz+rOY+uxTKrWZbx+L10tJsnSttt9rNPmNGg3x3WUWB+d6udMhthnGowVIUxejenq
uDb/sNsWWBNaQth1nckkm429DrG8OxuZq5wXyferlYdQmTL3CS+qgToMxc28FL4UsbVUlNUx1du/
83guu8Q/USFyJxwvhB1f0RzAUsrTusqQKh+g+LjG6ySxWlL6+EAEAocf381LPlwAUB14tKDgxqBG
gUeALWBRhSYLqQbRkEkWSd+vzrzJAovlAziVGnD5xaOKvnu8+o9VWr1cJF9LqH6VBAj0I0S6fkq3
SW4zdxCvujcRXTSp6hXJV6eBoKrmpGCbBB6Vek62Zkdzexg3Yq5n3vjN0tYr8X9rCQB0Qyv36tbN
s9NWn6CfmNeVnSM4qQhuPxrRyKsJiA76TIotlT1S2o/sF0o7KKMspT8vNkUzj/fwMxOZTdBp6zcg
mJ5lDE1lyVBnWdg9cKif1X6t0OfaQ85h7KeF4X4zgh9DTGo5aRfLBsSZjfldjXwKE5cs99vThKee
jlSvrpnIJi715rZkov8mGK48VAGJx8lgHhsInc3v6/zuhLbCPYfEYo8fjk5SN9o5ySNLL2FNKQOF
wdzgNyAnrtJWYSUmQx4qyPNhTaqO5VaF+rXmtQuEXeo2QAJGDxCXGOopFrFxx2INJuiR/iHfTAhT
PNL8p/yIQeKolt/pDwT9cWQct5Rz30JiSvowRVpnARm13cC9SPulzbt5y6ppdRgv9ikl8sO08v3A
NGguKO/czSE32mymZgCIweMK4cVxhjHvF9EyhYlyl8BPayhVLd+H+QM26Ly+Fc238Oq8hA6R+r7V
kJIaE+SvKh8MELMdUeaK1O4lvDkB0lFpiy/GI/+jkw+vP7fAqTLd4TLU1MhYrQ136lbnBylPlfDE
ipejt8MST9ssqQUw98WuiATJ91VzU4IZmLAVPgQWY6T5wQgfslqcuTsEZiNrmohUKY9E3hSQ0Hk0
S3ZSz6CEpjEkdejrXgbi2NNqdZbt/9O8T5MW+/8SQU3QGYaDUzvRY7MYJAHgLb/Ahs1gUNEjBCWA
FF3bzTJW+EbqI9LEGQnQmXsVG24rNGLGzjq2mvoQuzAHOKJz/g+EFHlP6y61r45Ilb2vsFfaKU4x
r72EWNNfQehoOfCVNs8F3qHUcd0yfEaPZrawDYl5hPGOwnYxVCW32+KCh06xNzQeh0RGVj7AqhoX
GASNjlj3iJA4TkB8/mtxIQ104Gg1qBRAMINr8TglCOi7SHdx7UETii793I+inq9DNGYwX7MNB4DG
GclDXeOF+DvLiD9esMDy2J1GrCllov2x/nWaHclCqV4N01N0bSFjK+n9vI8CFP48IOfwK0OZ12r0
SX5XQKbGzsuhAa/hjQlix1N9rfQCfXKRy55URdHB8Um8ZE3eT3iDzwQpYUMhXFDH3bTqk8dBtC/N
9Hl6uY6R88HP/JFgIUlwvNJEe2dYHffjzxaiIhpQ+zfdvW10X58L5Um3tmOSGa8uvn97fVM1Zgye
qMoGh7qRI0p2uOqNNdtxNmt0EswIBlVDzkYLsiRGYMHYMsmfvSJl2o5E8OlwM+OJ06Xox6O/ge2L
88xeiYiF/boflqucu1hAWEKFnVZcDKhpKiKepKiG0WeOu3IqfLAyj2+nApPlEvsHANT8JIYo2Q+L
/lx203VJSjzzwrk8YOIDgcTqWLTm8tpLjqPlvPS/DvySLIPhiJpdlYaavO1/e0+LLoTZVBN0MX4o
XDvh3MechKinaIBP3yYd2nEGxN3Ta9KGd+IOlEw6cz9F38CihZx5A9gnY5MGjK2qqw9smZqydR/4
LZeAiI4R87qT7xMFvq2BfiO3k3nMY0EQM563ETDh3c1fO7WLTmDDFaB723QWZJxxFtq4Fe+GKvZ6
A0MSVO6MgDwUTdU+l8HQbYAENCN6dGcN85zMCkhagZuGa1sM1Dz828YD0AsHomyRBQF2w5oRBEg1
jKCuEUpNIHMl+spkmg/BQKfa1qXzPjhpth90CpMbXLty2v2C4DPOqywB7w+PIuKiMe0AVGYs14Gz
L16yF8Pn9eocaC5TuabCMrxpFkVYVy9MwC5BaIbeFD+sERbMxTaGENezm+KrmGSPjT/W6Wrb5j+k
vcGNeC4ZpmQceV2kPDSPxTDe3T+xICgIp33yWbmn36Roo9qSTMf2E1hP5P6pB4313heANkgGCmwB
grxq5CLtPDpDTT3q1oCZ6Z6zCsPNCaHk9fE7CHV3j9t2r7IgsgJrVX6i11T5W//2vRGv85z/pm0y
BtROGvMEKMrVvTO3IwhfMpodkuFMPe5FYjpkJjFCl7IWnOzpeLlw4w5aUlKLjrEsEUQ/dBTXrr0y
m+ZRb+dPposcGm/FODkrFat8UZlPuTTr+YstKYVhJDqnCbxAOXJzbIH3CNVyKVjz07gTlo4OrZ+m
CUSFHgV/y8MdiSNNrsv5n2T8rV5iBHtMgb6eiunFNfpb5FNghI9FkksHrmWthpwvRa34faA9xs3B
Lysci82ziBBw5NWpFNUPqgDOUmqM0KpedFOr79WCM/vFZsDFNOXthMdXGIX036P8YFzReNrEn1WT
hv6bfOsRg2fTg/KTf/InSHvcBLg72p9q/g1omVW1DNeYqUSHw6kVNLOTS0piTWe0bCaGAk9ASVxb
NRPsiGSUaeGiCS7mp3oQYKCDf62FRlOXhrFapCENmMbRRftyzvWFBx3AISeqQg7NaFSa7ZQTU0Tz
/7NVJ4XDMOnr6Jr8i2odfCGYY//Gp9LcGDG5bvDIhODo/Sn7fa60bxqibf2OLEIssXWZFelIwDLv
ygPR4pGLsh26BheSeS0HQQb4dkLHgQazKYSdKud/Gwzk1gpEvFWyy3r9YZD4mcjfTIUy8oRKUII8
3Ftr9a0p3mvyhz1XeNRsZE+yckBSgUhFsEknk6ibr4qMSrYA2yBD9yxMEsSRwm9HakQr4MWswjQj
iYoXSOZcF6NY2w+yKN1r9AdifvDymxWEl24FTwI23L337SdQOr/QOn/3r+bf82OkVNJicmMEN9Cn
E0cjpEFgs93zTPycNEWj7zvzLPvWFts3p0x565qSsu4ftmPc37MOV9ohZjKO1/ZUYqAh22vs9XJP
YWFhBkSBCvaseaSSjAj3X6SzHu6NKVsV8ZdhCuT1bbSBVfT+s8f9I7hUIh8uMylrvaGYE+prX9FM
ksJFwI607R913YmQxCpYCGD3eeDEoXMXssg7yVAjeflVXGuzsBDHUhKYbATLj4r7ak5I2TmwHUOq
ySQcDviQ5t3dNa7BZciB6y35DT5+gaZ+HuprTENVUgj4RoEujYeUXjnYfom/8OWa0aWDVekmS05V
KCPjsA+YnDCG1X0EfViscVshQtt4yYLRMBAnJIyccpgwyQSTAzAZCe6ymmWP90nqnJD7tODrIz3I
uN6rqd2YwA8+FEcT5XOBPLyQu6hVbM/kkQZFGwhsOHJ6N/z6h6jZRTkE09oMq3kjhrR2wovZXPlO
SuYg4G0AmLMQxs+qa8dampBOl9LmoO7rSj0mWcE/tmaSy7vveC4MDRugeWxKPl7nmHOL2izhFp8J
K2JC7JaV93JUmGV2HvPkw468kdLzAYl3oXKNbO0M0Zti5MCzgxEUCSKkv0XDP7iorlGukhVXD9ap
ycBu0WojCVmhenAujDgcTwLHhylVk/qVtLDWdLvEuA1sw3WJz/D16JftnICYBR3i6LWXIxl25NEx
UX8fSShkiy1i1Apyi5X7Ue0TDfO/3ORwwFn0OaKqoo4ngYlHt9GeTdACiZEm9Dj64YcUmqq2VJRF
Zv/IKC81Jf8nknKQEXyCQzp+GFGzXh/WFFSNbTAT8Z0B45/FrfQQrlZ6GNGCIt53pX1dWl5eYQ+C
ksrvfa6h0/MVPSRdnJiYOajk6n1u6h2JERXwXLY1/cp43Yrez+kr4g342NQQzh9exK+4kOEVj85E
7kU/5e1yIqPMNN/GNgdBRgsSBjoyGifyPyedEZT3VTxmnVdlTeqSnnVCRKTNureNjTqZsOnfSyRy
ZmOWMYaXJwW+APwhpayezg+9nv0w25v7TedCuya8/ONE+gNWerpymE/kjDrx9I/UvjZ+I1sbYybK
1kqPuw3pQKkbk/AzylfScwJj3D4GnqdWChGN/quri53uEt6YRxDnRSDXL12KeOxH1L45CL3jUY3w
He+9szjK+ZWoEdwGWtCTIZFnNZ2jFy+bJ0w+wIAzWOVrA9TMyIcnM9BZGgLeJaKjn8cmvP3eaFPR
DKJZRwmEtvizrEvYhZCuAqlBHCrjNyy0SVbNHXy9E03VdfyF/QzLXc1OuoBy4l42McRl7mgRCDUe
iiiN8XSiZApQAgyZS6q3LkymKHoQYiqskCNZ5mGw0b12PXtXCQ0xCgC/D7g1yYChmP8UXRlqw4ul
hKniBFpd7FJVax1eXDpojLyzZSXlvPDY0ZWr6IQhEVPlrrtx08N0gpyNyCeVdFDl2ZM815BkRzQ9
0hwil0uYG3+Kin+X3jpoivAPIJ8qdgkE/npeFPPft05D58z1gxpSqxBvmH8R5g5gI4EpzBq/bO7p
Xx//XZfiMBfiSekg23PhcLNgOjthJPv6+PXCCQ2rTvOjAKarygHO9K9KDiCoPkzFMelpkE2KzYx9
V7itVeA2dhTLBWYpJITskmDa1ISJ/7n6MwKZyLR4oB5YB0fH5P3pKkq1lAp9YrnMjfSi7l+Musyd
6jsjYjC3b99yOv6PbcRAXVFocidafNAoS4HgcdentwbJ6wtMS3rbJWZhCaJDXXgCnolEO544hk+c
74kh+gj5ZyzeGr7djrFcC8IiCpacckWbi6zrH+7CZLkrs/uKf1B2eJgcZYrW0VyUjj51Tr5gfLYx
xwsUOlzQkTMoSxPzQ+P45dWCk4PspPcJksUx2Mmif/bG5drwLoV5HcVv8eQKsgkAzb4aajKDdia+
A+9DYFMskQqnZg1HWepjj9AP1vxKvRhp3lcP07KA3deK1mv2aOV1t5R/yemCj3dd/LQiQw3twN7t
b+reFM0fIUiyCKyTdAMqFEt4tl3FUWDmoIh+WDpqpURB6Vu0h5x4WtSf2quvv6nhkGoHJ0HS2SLZ
+K7c3JgLhaAzn08RVmHWZ0eMogBcCCy/F6g0SBr5taVnMlYPN80qqsTP4p5cuGEcTMU5gEm4iaBq
1XF1+xtKhQ9SBG+YGzqbXogZ8yqi10QO5QUaVZs7zIIQtfeEgXWadKv7vWe8JNi8z2AhZBHBPwMC
hB+F9o3ByGMsviSmXdj84PhVUwFAkXDL6TH8uhq8xudFggWkwukp61FUx+4c+7XK5X0yxEwXnogR
/Hcp+66fC1TkkUj5oL+b2DSoVhqhc+0dazfwYrByoUd9Lz5YmKQLET7CaiJNii9huFqji4w6+XNZ
2mDI6ZXslqs0kf09VoxfotHKXPBmv12E5gKnJ044KgKtsT3Wwj7agcDt2G66yBGfHUaHIZ8vTB8j
KRfNPb1PXmDPohKYojI6IOoUjFzhKeMCHSD/P7TcnqWLVbFgTeYSiMSUWWJdfGu6pFpBNtqBoM0m
F3VjXE5krb5csU7R0hRZFek9UKhR7MDQVCLcpEO1sfLbzk+a8Mlj+fJA8MmIFu9kka+1lU/5UBXj
QDZWLsYDSTHKSGr1ChBGD5OQY4VIW7FdRPW4cXaMX/ugOrL6Od5Lz7k32lokqVczr0bcs4imnsrS
Nh15mM5wVjap9DNiJOHOCm8VNjrs45OdDxbwprHHupklRbm/DJUToHzuo8V2PRM9fU77Mhth7cR2
TVsJtT/Z3/doPRbeJ/BnOXHY4wqFXtfgve3uBlbVr1CzLMWFU2p/V3tI/9hYYcXm71rZ7yFqczR/
bQdxUFs62hdcAX+mkr2lqBXIFktc4DnSBPe8hm9EybwX/JWWPzs7dBlNGv+myZqayBC93IhRXUYC
iiQ1D4gR0vVg4B0HtxbuEqgyvurT+DWFnCNY75lXSPHXXxcod2NHPf+0Sn/I95jf6L4NBoHBudIC
qmgaCXkLALIcRgHJo3FiWH3DXOhQECwuJ34sw1yLD8iHEKCOjaKp8QaAQYKfKLNuKObKF42zWcgY
8jhs+91Kp9rxQ1AT+hQLeZFSWf5iaZI5VVvbn3kmDxFvuff18HgL6jpf6MNnOb7UaRlh8CA6fxor
Q2/1672NgIAvcXWddUXusxVPISHzRcvOtVQglOc+rWYsuY6L/0i4lXS65bP9yjH8bhRAUbt0mIcL
U7/YMsNSr4jaPRfzhBpH5QDKihMOTWl716JhMhxV2ZWk8OlYvWbsTQ0Dg+3ht3KdP6BMywU1yQJs
ymKEhRbGkmrwg9ycaW5N1y0vdgXwGAO95MlcdIETLb3WxBCgKgmg7btDWhrBIOXbihHxPGv1xoi2
URCRYynUjSCrdsOnR6mWQKDTblNg0T2KVvH7Kn1weMFHHQ30Y5fEOMIdrz/fsLMbJmwDzxR+GS2y
Y88pw1pPdJ+JVpE1pWPYUFABXXe6kAeXoaGA5CwFDm8n0eVg+aldYTzn+hiohtcUP4bhh821M1LR
yQZBNTQ5wqueLRGvgGUh8A1Zc+6mONV+fsn6UTe2ik6X/c21hs4m5MAC9tScmz+EwfnO2g5B7FCb
nzDmyU8uly6k9gdL9IfibscsrWWxyTwHPh25GtzTtifjXtsvMVNFHanDNn56t0WOmViCqaedXklz
DxV67MmfS4FJ46wJgd3csgCSdt7M3L9S3umzICTK5N72KbsO2Uua9aaFXMNOkzKNIaxxj52oh5Hu
pFXMcZsmgyDJtolPT2JmpFtj/lnaV2FwoaSFh4nssSglJAs8U/SZ1KePoFGXAkoxyBz6NqLu/5Pm
PQ/mm1PG/Nx4zA0MA6JT0tdhXf7KqswS4SfKNYXFPjHXA00JCs15tnwQJfRA2tAJKAq2mAJv5iRF
ian5Sx9yc5EupE5VSqQ40VqTzuOGXe6WK2pt8KPSg42JuA2/KQcrqj8WP4+T6BSVQypNefxznBPU
CeEbI7T4g3zLWNkjuSEn4amk8VfylPOlqDqjfmjQ9m6nzI4ug2tfgdwgWgJPqT82tnDsN64hz0te
OQcxTmoQgScZBX9Rlwoj2lT0SqTymrQ/s6MJsGoLn8AZA8oNZbKNIUQiHdhnAn9oMccAhEOnYsca
7snWRRp2ZWZaeiS6KFV6fjNbGFd+c1q1kXuXYY2+REf1HdzmmQiO2WXR5LAEN/0tYzzoOVORfCs0
LgiOvvaSsSzm9STCiLvhJP04ql3ZVnxHhPF/knYmlK+MyQyDtDL/0KmvSILYEEJ/8Gdm+IJCYFtQ
sINR+z8r3jPRqWQW1YVlZ1RJBJOdRXApjkKDGhuB7MS8f+n9zBYy9j16nZOO2GqZioXeA4s8MC+s
CF32peJwwOB1RGbQJZcB9BAq9RoMB1hf+i0DadaUc4mO//ez1xXEf6RS5cNN/5EBxNhQK8lwS4JM
jqeJE8s/z4GT7zqpQPFyca6b8EGJW+V7G3VVPIt2aXCynfPXIzspGgy4WJjtuclswxM7gJoNbKVV
rjSxqKuAaqgbEybEcTRFIb5DnBuM6hQymC15jPiGIBVUQLTEstOM1tYGh0+NZXPDT/BshAAkchSN
hBgl9W1aHtxuwbrhJOQ9Umr9tQpwtQ+bzcSir+dhuEsHko1moSjGTrMr/XZ8Y5o0yOh9bM/0NupR
3Rz4fuL5zzSSLgwdthotDjJqNhCAgnhIXJ1YaL0IIDoZpuaqU7BNgS0y3XbINElItngsqLJy3GBD
bnJYIFl7bO3iuLBfLZI6Pvut/BPnutBjoF0dLrArvu5/cpCBvJTDOHukKElWpQjAwX14oJ/3HxLE
xzUkHAgAgqpMwyNP429GdZ2zan5NNOvFmrQLk8dgJSAKM2XLOKLvm2pZTODxJqeK3HQMtukZ7Djo
5gYa03R3mKthQ5gYVjFRWKbpYyv7MvoSRM/jtTjZzAPPQD9FlaEo4TN7zZouJbnElFibX4sUhY9g
u3jUC1myJeIrl4BvYQnPdhKVXXgyLa4LT9e4d7Ik1ekjDbyKGxiZ/gpf+UZU+4VC5sbLurmkzh5m
QTEvBqGjjDY8ZaePrrVTFn2iCgInIDOvfTi5WoUxM1+PLqnQaBUQ6HyesR9VGQEoKTrKpbr9qbp/
Yam2Sp9eYuJr5qBdMU/hvyT60Epze7jmDWLNq5eZ+mBwSU/xIQkhd8/R0e/aqivt0F479QTJBiFz
lEKtjqAy5fwj5sPI8k/lNN9PjGbxHR5mgAryJerWmOY6XwZ2Xk9EWEt00CZQDs4Mxj+/qQnqACQL
ZA0FzTcUHHPE86ncjri9mEynPhLKjyn2VkE4oWmkLF24LVffV/6YAgzEQ2BIbJ2F19ctH3UnD+Cs
hfbgETwONgzpzQNZ8NOqUHFq/sc0lQo43QcP75c2v21z0DD3t/nbQjpqKjOTCKxvyvEs+Krigxjm
GvW6/c+UaaPgiddWDwhaOwVNs3ov+ZiT0cHIppNWgV22bqb0jGUwcEdFhy7Ka7K6qtr0scIaG1VQ
RCdSzriYkEYkFn0YGFngBKwLx/p2Wb7P92TVEeDY7hO45eEER/YfytZVZH/Qn47EG97h+zHYFpRw
B4ZArltxzVnJmrlIXeaJjrbq6gKL67EpDGWorUmyY2R+oOB94ktjKyu7h/6++b0SHUQwP4O6MEJ6
z9hCixKYRsmXFOJ3BmEO0sVtQgqTwd6Fxfx1r5mi2JpjxVTBQ/HQ1EDPfEF7FN5dd7fxiSVZVMB8
HHr6dfcCEX6tOqWqL81Tv0dw6RL5AK44w+B7FeaEYSvxkEC1cAsQf4oPkza8efFA6tgl9JD23+yq
uluxokSphHKvHXXmmISGt1E8kAtBSZlDVUrmzhkpzohdmdD2n57EWkMkQydaabwNwLaFp39bwZMp
Lr42JFpAmktm5THR/8fylsX7JRwqFEZklfivMjEb5uGMvV3RfQDCVjXLdV4fkAW/RcuakPFp6ON/
uRF6XyyNpfqm/+82ugcMq8fPC/S0DRp4ri/+sFxxvAkSXJoAmUDW7P97f7ammhuklFmkCHAi97SJ
XBDgTX/gexD5K/FGwo9LWubjL15gfYedU0XrC+fEjtXB8aUJpcnevLDvOL5qaBFN45TFyQ/qmFqI
cCx2eG3kK4eS0M23vvZk+8Pcls3qbL9CpyCpY2bbSbzbxtljsa3oxt8EHWvcC+wvlyULKWFmYhBh
Y4esIsONFHkh/1o7UOkV+lGxnZotU5LeFHykOFnQKMMsy2icECyqqBe1GOCIATinzb5TUG0OIVEX
OV3872GACJOO4/0b0qc7UWgQfRLSgh/Ca6/Ux5R6nhSgVP0d7Xyval/YAI/NfUk6tZ5VoG12XuzD
Kq/H0cOGg51QQu4SiM9L+7qzwaPDnXAn3TzmGZJIr7dfGrugFTmt21EIWAh0ZM+TALgtBwsLT+VV
J1dydY1HcKFYvJG68877Yctyso0sWf+vD6lHSbPr8oMAWiLNqJqB8nmZmXQKA2DvTNMSA8bY8i1q
t+nI4K7aiSujrPYHloV+ucOW0CWpTZVQzthdZdjAFWKQLZluJ4b4dzUQjwQ1as3LHmN0vyMRFBGE
iEyhm7myp6Fr6MZBOxp1qMlmoPjaxy/TLIS0N0nCmL/9bDLWR5x3FblDXB5Y1ksA5gnFVy/tH3Zu
xiRyOX6fsLjxIal0tK6jGyVF7mj0oYdMRIojW6FoRUgMBPJJVt5WmOYKWFsoiG1MrxYmwbKtpg0A
RlHpgcgzbm4eWFqtrjDVOnhyqDEuLcuSWA9DPXAnzVW1Z4SH1zF1iXu8vJ+B+wzkVzZyzBzYN/tM
y9UPOEFsTcG84PIR0uVQhSJAAf9XqmyVuAVjNzwE5F3q9lqRnK2Y1oKsjfeWe5UIHcj8Bnix+po8
W9u/E5PolQSrSS4Wvyo8Sm0UCPVOPy87DyxCRPacOYWXBYW/X/0QJo5TdkrVBA/8yYcV0QhOZggY
HOPGb3lo8poF3kc9OGhSwSn9bOe736TQP+fJ+Xvs5SZaS/9kTHhnB1YWYHtei6iLlzgi/R+wzbjw
8wTc8Y0IcnO2PN8BySfn6taanM7tqBw/XsnQhYwtppBR3zhg3XVWiJdbFjetleXuiA6wVyj1CKM4
xswgzSN/OHV8Blz0pwnPn4cIIVrAOeNyx12iJpWO4mtIPITS/SlqUckuMfr3VnWX3rumHmOZ0SjT
cp1i6z1AgCnYqvj5MxzG4xhxSrJecvPECyNlhqTvRR0ZH+vbZg4riDUb0GHxLNBoZCT93YcC+lmu
vziV4Mlunk0LIpslfvaGz9v5qpPKoAVw/d0diiqsI27Xd2i54U2aznhevrDNW3zIUGGGGEHHW7BP
WiHC/89HBggLodurwrx8J3DYM3Q/xO/gZnAd7FMhmXMD+SKjMsCbQvInaIPFgLoGrsSJy/JAvcnT
Bprq8DVAN9QxGBxIVXGkHWqSsPjn0gisoY0YZ9i+mn5jKlY8Hxn6lpcEmQvxVlKjf9MSi/hQmjmn
zxzBpIg68TjLnSQ0IFCJBO6oqeES7VzD5h2qW9SD9jh9hxY/Nf+RjaziNQ0URwcH1d+Kiad22aH0
asmwjml5S5JUFWaoE2tbro8PDjcCBegAHbw+4VL3YQYfyyBHJOymZSRLUj/HayuZD8BYbf++zbN9
J9lI3rcnj8FFcPQ/0nlhB+uy1QLixzkAqsBrj/SJ1Uc6Yv472Wh96F+Ow2CuVOm7IywITqLwiuMQ
E36rLrM4kD5REWKe82pY4dvJDq3wsaaylP0NW1OewwA+4ygYoQtXE6uE6kD2T9PmmwLT/XYX8HwQ
cFMpRT4f8SUWNSaJwRspw24lqBkQMpVuYNZaWC7qBA0VC6Oq77xcB4GSpJxslofdA2U9AGZs6iBO
NOzTxn/SJ8JVLIi0fY4w25wRN1UCSbttptxd7dj4lxrSPd06YYzco6cM/25252vYAFlb+5qmHDZS
fiK3+L/JXj9UNuZJmcRPn7GaMGdEvA/d0xqFHdy5FqN4PvH/iMN81mQILi0VaD3Fa9ervi7Oa69g
zv4bvMKc/pQbfUxoo+G5jCM4O64Sj4j1OO02Mj+9AV/ucg/aIhoM5ZEB8P0OrpMyZWlyw+emcGg3
yfUBgyAtJt/MNi2Dvufn+WpErOdyc18o2tr4BNU54BNxK5BRwgjeNmy1Dw8TlepCQ09tiFQw6myS
SryfEbdZG2Cyp2laAeLbohs+1CYgmjEfpHLblJwexherq9TSIJFx5gD7k/Ec1OjwuoEf+ePMqFj6
Ta3p8zbohwfq784JrLiy2Csyw/tdD0dsFjZzEcKQb9MSWOVrFwEepPn1D0Za66Kwu3Zr9S87XwHB
kHmaCsnkgp4cyPISAAZtvu0b0/elF7sSXKOJhbn8NPiTMmtQaiMbOiReCa5/8NjtdbTxeTwn6A6a
0Mf/j0GWVDKXyYLAqfq4YtBw/YMqFepgOwnlpUFEXFfS0Ub7IoJWKcJlyl5NYw/9byD5zvlpr18V
Izqdr4tUS4S2c6Oq5jvWBToj52M2bx++8lrigadmMQ5eZXGcANfD3L67E4SIeI+WyVist8u3AAou
tsXjvtcM9k4dxce5+JCHOxdPJu19DXjSKs9IsO2FtIKU+kpACGzBArIyd3eRURXmwE+w4hWIsR3i
QDigNDR/neD2DE9KoFhaF+NusWLzSbRYe6Pcf8LytntIYnCn7lig3wk/m4/VZcGrxTHrKfswaC2P
ASxG0K5G2qatESe7Ot5IQhpZG05A0XeewgAKrbnlUBxCT58jsDYk//bdYmBY6DOrBN1NhNSpICT7
wC49HNhGkdGBXxmqhDrQoGrEqEJ3LuV/BrCdy5BCULWIpStEHo0PVelUiOPnOOM4lS/hvh4dfTXl
vAJVrOVz8RPOyVZBav8TaiCWx6T3XuRdu9mihkmMhA5JnBXxKW0AJMLAJt76h4PITfS12wKDZGtQ
Vi68aWKr7oDuff3kEr1sm7RC0kiNkVVKs8rL0146aeof/fGd67vu8vxvxq4e7hTI8gbR5B0RMT1T
r4X5anZPhMlgWP2PCfCALgKJXeSCr0qVCE/cAFauuY1bhu5Pcd3Khr52lZ/KEQ/pCFk05OeBSMiA
ZI3qj7IZikrEydsFPsBOGmsGDrL3+UWUZWctUvGDWm62NPt7CJeDlZ4R1HldfoCkof1ppec0Ixej
sZlS25BUO98/CJsIlNU5AG+2UAX0/uYk7/XzfqHdtDqNntQbymQge0sJj7Qfn8tZZFNcuoFbJuoc
etaS7UbC+IbGhJqceOpVGhuoJ1qJRH/94Mv0e+S63D68X8Mk7xWD1cMpx5DhCj+c9tQlNAkj56iV
OZVCgtjpLpjU6tiwh3+h69R0cRCSxNa9ul8+9SzjnUB59hyui1klw1cxQMDJtyBhJMeBS9aimKO9
WZVnddiLd9bEeN2H/tsfBkmOVtC8W9G8+Zjx+RF8OlrSL/dxNhlsoVTOT46rhQ6c3n1BwkrEHKO0
S8kAVrPFDD71mFPikkhdplkSv1+4GhVNvC7uUOS8QD7GlF0fE75dcX9xzDZ7MoBLuIKcX2oevps8
c8vlp8xKOKa6xhg4ykmzKlhj/smOnqQfYyBube7oCT7u4HAwiAnna26Z7hDQMa26F/VheSVwurAA
Xwd78x6XHfOHJzXM4ZkQGBJBlgHFbHcbjbK7n5U9oycaN/0EFdezwKV1CCaK9dVIA+nno+Z4BJSo
VIWu60VrWBDmQkIL/8UsPQS6tM1Qa+cGDmHrU5IsfupqD87uaSbeNd5aoMuUjdwxSaRYFp4CUgSf
p2Y+r5k08oDZCnVFp2Ur2Tmrb8Wlpegrl7gCUGQsd4ZkypJ4o/lXxE/AgLctBYXhsavSipibReOR
NLm000BjGwcajWmuDbYE6oGbplI/eYxFPuvTG9N6ANXoF3vHonsHv8S6ytzK/0eg++7rPJOOSw8+
lHms7n3PaHRXcXyK+LFUrDer10t2ilQ+utKUUSPwUCp1Cu4CoG4dcp651Zdocai6L4ozsSzHPu3H
Smj4IKJ5TxxzTbB4/TVl0PQVfqtMDMGtpoSnc18ouTv23CBPe5LDPH1HV21Dcf2elK/nhr3wXs32
VfPScy8xg/ipjFJKnJhTMytHSRcyLPYhYNxT+L7tY5+vpy3E8zsLk4t7UeUewY3Ht93cXrJBOwd6
srXzN8fLuJNeDdVBDXYZrfZynwqVs92tT6xhqNxe7lhmWLF/7sUBKb9KU9iX3lGa5v+yj3tSUKK/
1jHXDj8Zy/FvT0ls3wlyULWp2BlYz4Fv5W1yEPLVCMWDBj/nGKDU5wv/Mv3B500pl7zg2S3S8ttZ
lABrfrgK6rBiWbLcage8KwLispGxPaHbnKeJAibqJcn5bd9t9BEhyPBfy7Rj0qGcHzEAybVatlNf
jmKvDbVLDDLz+YPtaOAp0QYCYSAFVdHKFcuaBa9lBs9RR0ZYtAmvL0Dqi7GtNPqsOee67Xr70diX
/StrYAUmoxlzqAexYy0vjYpnd+SQ4GnO4yNffNZT9hIdDLYL9BVuYzIFZVNcrnSL2ajHsvVWYWqd
DrQ4EVPYQb3bze1aZPEsWRVnF26E0GhEVFM97IkWJHkqYpnMkWEr2q2YdH5hWBbAlcf1y/IeQbpP
LsD9d4o+z/26TIuhG9MFLnCjCLRwxHkqMllrp4sQUR8M6vYstaWTO6/Gc0w6eUZp3Qf/FSLPhh0C
pKGJNQ6Z5fy699Rnn+Mb88/rwzhOYxpi6NcI30jAQTABm+IgquaOGpmykoUTYJ9rCwYZ7eYlT12i
UL71QD3sFMDxurs2H4P45XwlWVyYH7RUdLIDj8lB+sLGYO+Vk7Q21tvyehUND+O8nG0ne8PNBQMJ
6hW3mlndtFidWPaTmQe4nlqyxfc6J+mV57++YAEzMSol7Gs3uW9Ei4gLUVotc+UQQqXIWqxaq3qh
VHR6hNFzP71ZYTt4oF+HepctjjE58G8LWBYyv7GMqq3C+cjWmR6ACqOB0oYf1BwwVtXa9O9CtV0X
v4ks0V83dJAEEpulw7mpLiKbW4UPYah4X+uvh0y2E93C0GEFU8EpH6si3wWow+H7ZP17A8FdzZYh
JCYe/4ZOQSZORyRTYKynHnxXIZXJ1TLzW1ozF3f4WEZuKI3LwsqFVyDgc9NEYcL4Nu1Sr9qavWLl
J8oObkgci9nTbroAc3z2Y+4t+7HC+6iid58kKbwo3CnToH0Le5uBIiINLv5+4J8DMtlGVl/F7KTk
MbwGOi0NI8TFwntOwX5yr+vW+urWQq3m68UiH+7nLvyAQOY+GzilZlArU6RJHfSprvZHfk4ioHEw
+umNHqoC0bCB1+zt3eBZfy0nH5L2bN0/nq5xOmnV9EIK86VP4E6h2I+g1SPGOykRauowJJqa0yoo
SY2OS49TPGjdESiWFDPTvb53dG5XrNM8mTlXWGn+it5GdnxIzX7MiQUex4QZrikHUQINNCje8GBl
inVwj0OZZwCM2f7f15VaywNgQIfB7wtl8tyRR6UPQ9wOCDnI8MJlWWPAQ034FT/wgDiPnwMGdsvp
boXJSNLF4rVwSOjJUavsd6IT7j9m+ZenNfEY+nnyRdX1B36NLHFta94HqNP467mBPVMgsmdEZCCg
7j/bQzZcSXiKMBbnagDI3hc5a3au4YW7yz9YMFYyykhb2TnXj1NIGLRGq614tlaMGUymhwYkPrVK
doTLb8u7AlObGGLm2KEKDGMQqQ81BapGxR75cLi0SnYJK0NTrQtmkaJA5pASIhvjN13u7pjiHs4Q
qiPaUNVokd8fGo6r/fjCAJenDDaULzBVFTTUkpLinJTma693mx6xk0fDIU+UH9IF5RsdX45rtiiP
PpzQHTkAiVWS2JvDZkK9cjx0Qx8F6hBr9Rinrvbl/HeMpTCfZatgl1+mbVuPeQXF0ZI0RVLFx0x1
8XQxsjbEh1nnVQG9anzbmHg4P6BEmwlFRx7vXcfxt9ofl7OmMYbcOQFbu5r+6EyDbPUdOEYAw4TH
2VykL3JfUBwvuQpzkghxw043AT5Z4TxlOVtNFa3gPjufmPqztqJ2S5cBrlOEJDvtZbEApuFYDoWw
n43NbCs3cmCuQSi3OtORIAS/6ZYWWHc4VJrwuue3Niipc/96voSdDtZjy0DzWUtFydXoNtT2WB4w
IErCfi9xoxFlZQEvMeFJ3TpTFpnQ3MZJk2iitCCCnTYXLYCtnzsWXNe6OLrOHXQbue9XiCUq7izg
b99m1cVFhLekShWCRISUH18LNgyom23PsCFh5GIgdrxsBphs7R2Zw889evztGGJ2KVOCaguPKE43
LoxBO499eSVGQG01EatXee8QcV1gmUuACQZrpvBI9eZOh+8XI2NDSxSdz2qiySt3R8qA7qbiKDaj
gUqpEr5hSuRLAo+Rbnhf+dVk/3Z4G21+iOt2WPK4KinBx/vNftF6pnfab0knIvjSUTY7zI9/nl3x
2x28zQzPj2SlP/KdP1zz9raVG5uDnMR6bn4tx5dLui+0xU16VNxn1sorcI1FrwILvjGhtGuTyUGt
4Y1uID6wXQZhekEJmIUKNpjybC2DwgQ24yxht73bg6mbclFgbx5iUt1hZV9rbXOieb3pAXHjvkyk
9C5Q2w63OePuzxCN/HwtnIdQI4dCtQZB6d7eCKqFrL7cPwKWIQQQCeaHyIjHLMS2PSGU5AAqBp07
SwLbkEF4Uno+ktPMCquAEPyRantGcAlUg1mVYXhdaWKR4L+2uPZUHd/RA57nFbHLRjJ4+kNUKmne
oVhTflvWK/EwWEBMbShi1dh5ikwiczmw4BARyKTWa9iXUScp2why5E8aMcS6FjeyWnYL8DNB8h9t
hm5jn5RyUe6nR0c239JEDReUDYPEHgiHkBigoq50TAXd1JiF4EipPzBqjw+N/ld2Nm3J96S+rGy9
GdhKNq+o7FyP+aLWr9N8knqTIbcwgnaPzXHzEzAsrLIEIgrHCmcM4XE1AIJkYhTckdbeTZZZBHHt
4IpOJ8mL7sMXoswK4JTC5d9M8CYd7DSkDN3MnoW0JTkPfPJkiZRnQKUan/6Od5AeS3XsaEBGBwq0
Pok2tf3bD4WPriuMF3gRng7hWpTWxthwix4hEwMMtXjdsaNqcs7F417vBXEuDWkCNoSBryalKJPh
K54lDg413yIf24LKdF++3oPnPVvnB2C/Fb9QrHRkXaKH9V2Lo7S3N+9qbSfZEz6x+UGAOa3A7ng9
v4DROSPOA0kyA36xTrla8/63qu3xSuxWjlQ3w3K3zxCmeaBZfbPcx2v5cSNsswNZdIzZ1jK6+jRM
DMoDMTxuS9sd/KCVIjbNPf/1qcyAqBbrsUshCuf6Fx674sMku/dzNgl+07j4Am9OH83LDaja/tAK
FefUIWHhMPK8MSeYOnWR24gyNeqRmYecPqDCQlVHSa4tV9eWt/laGV384q2jdRcK25X3VbprH8FK
im4ForxHK+7qPyuJ9F9HLRFbVvCsHzg2d2CjYFwNcr77KICnrVMKUJjpjeZCmy/STvt1mUbI5RCN
VZe/0vs4CfH8OBq+/tCVZowuFrE5Gbx1SpUaHnkZN+gqpsVesZpjZsr37jdf/qZNdwaR5Nl4FOAg
SK4px1a5Pg8VMKi1sls6ConePsK6WN3sdhfipcTCaX/0YAPcFQ4m2+9e5xe37TQvttpVoWUFZbTT
d0pU8I78U7YrUaAmnAaoamsORVRSQRyPVQqdjltp/Xcll9vc9OgCNgpPCN+TFSx/lPc485nTRkJI
kjk4w4LNTgCRE6PFZMPu+tfMxBfooswYVMhc4i+EUgI2DhG60UQgkL4vGv1vqjQC/XWk0AZ+r1OE
WJwil4Di0/C1GzPn2cwVy5SunApZ1n0rwQQRSWKh9al5mUOb3UW1S7IxTaoeHpXeXPGoq1sZhOk1
EIO7uR2Fq73kGlPM+LKQP9ocDKckzWaQeALyolSfv2CNB0NgCPqlsvpQ+E0chS6hbFIebk+Lfzj4
2D1Z9OEo82ce8kowxhxq0Kvh0E2u7Ty8ypDWDYzv7Yh6lFV5Goj6HbPNv01SDW26VnhHBOBKOXdy
H+SGzXAJ3mIYA3i40vBn+OyTCS3FVMhLy0riKDozJVpYNR6xBgDUjIgQJqTOMNF2ZN9GkiK/STQp
pdIkxMHVcgAJ6HZfXnCOae4eLc1tzIlYQxuY3C/owfxnR1TkzSoyoAO9WI4vHN8eByJ26Qu+cY1d
XLBOUixEQ8ompmuhBtCa44l5BDF7DU4iDFuA+2xRuIwLZ/9f3sBjzh6pATWh+TRqPuXgtD16FwD3
rOXwznnrhBVpGFU+ALaN/gLqaL5Oi8T4I7v/DjJ56kVJAX6Mqx/UTtjioe8Z2v0Lwt8BvAIr5mD9
DSQmDWPRugpgr1N6Ht9mMMGEnmwEr1ahXO3pL4BD74+Buw+qEsUDYwvZq+rk0qlaP8TglSpJSCna
Lb0tZTFWnSmWGmQohPsXsAzuvP+9WDcsw7Ixah0ujiUF3CWGSvqJkYe4329D+B3HGASahAgC+42I
DR88yL+/EMg5CCErRl+2U2OwL1581DnWEi947yErX0/Ryq2fgK3lXKyAJ3IvgRJeuSzknpWnu4Oi
DxHoyneCivMERA/4tAfDXt8C/I7YvN/TsgJ51juN1mI7aHT6ME7g/osKOPVRVg+DaK7l7bp+vNEd
CH6o2OKX7CH3MjghdqyuwDIgFLjbB5RyffVDLfausDj7ufNOsAlwPEZRV/wDnJ3q2NwcBRuJl62H
4RJJlFHl1kmON3fHlWcfTZOl6OKZmkK86oZWhxAT0KWcyHiOhKuzVhgxP59VVbqF9EE3J5sdNUaz
zn8LunEm0gsr9TPooVc4+BhtP4MvOF69oMcRNNWEfe9p2AL69slt0Lydxrtik0aHV9ZT/FxJ4Fb0
u+ahmrA9q2P1sOlzz6HbkYZ0NqZynRapEP+H/OoOgA74pTy0oATGO4T7kZonZDs4Jqx38Of1I3tK
XKaruyQ2qhVXO8g7cBY5362kWCLmGsUsS8MmlNcKjeoEqgYVuUlSeEwDtGsXmH1/yrVOTXFYlLr/
Xpobi3cVf0MMN7aozxh9vQpwOZrn9OyI2lL4E+dDTIXvYSdMaPoUfqZGdlyk7Ye/s2VPf5VaqtaH
dqHKGtyCL6oSJ98HXU6Zl5TuFgzTQNKH76N1tw/as6rdAp0TgXzuzTp3aqokKgcwoGsD+RipdxOw
O1gG4kQbZmGMYWy0Tm4tGbgZg6qnfpF1yOZGWQiW3oAVHwwhFarQsBDKctp/jbWXKgKxjvMzC5cG
C6joUs/hgUQNVVkOzIU/G4rHL/KEbO5O/bi1R5nnot2ExNSwuEEQ1Bx6lpNGZBDgdtBh4wQHxpvj
I7SIlkipscsRNGKRZCrZfKEBMZhCmSLYAJjY6gOQz++jNr979iIYO/A6NAcLJDUrezvranh/LPSQ
zp/EonYFVuWtLt027UpMr879oJ0KBEpWr3T0YLtq14g9wMZB7vdIm1hZx2rLTuQNcLPkOeV3shrs
fxMfYQP18y0ehSfuN/III54eF15BxqXkMx3//w/331zFtJgfRnrZs/SuKI/fiHENsHufMhj4v3CH
K1oI6enhntUXsjkjBOVsBa8pnGENV5I0X/rC0uTCs+pFsOCy7oIatagAa+llb5NeAcFJeV2LhbVe
p/501DXKRGFuMPnN4tyG8PpTX2K9apLmvnDh8TaDpQwF1jW30NNZ6Uo4yICQmvC4xlxcbZetuCrX
nWekb51VwNMUs7urKs+LVC2cmGHVsRDETOetCePb1ks6MncGh0QONpckyyykOVuk0vIBZ2lzLtS0
nPUes4MUXF5hY2AtwKzMvEbVD1cK1ZkhflFpWKD1ExtTfvrQ4+cdyAzt0cZ2EmsoUPTtu5FjiQQ/
l4OBttyKHr6PceLaQuXH/B8rAC8chHbWyB+g5JpZQm6C4u52gkg7zlSarl4ZSNP6ra5W7F1Ey5tq
y/N4TSoTMUujRXytc52JA+o8pDi4sVGxomihGcJRVKMkUds+IAtq+KQCg4BXvIR5Ia4skiCy+00m
TntlGURNpoqQLLCE8hXZRr6RjPksJM9w6xun1uAmitKHAtoSOgEZFK1NgVg2WjHa+aXq/DtYkOnI
O8dEjDHz2Dov+8VUqan7fLrJylgwtDNPwwmveLIXdf6a8qJJKJhJWxNkZnRj84IPmkpyThA91BXa
/KRKZ8SyL/Yps82qN0B/QjBkB7xx82tU/zLWhtjtcRI5ZWLwBOs8LmPeAfRpfch4ajORBPgu+U+V
irEPh48pK7a5g3EdF2BR22nfNH1W0ay6JItV6lhyB5yt2L7NgS2VKXWnCZDjamlkz3fRE5M5FbEb
1p8ppg2lMZpTFKZt6twqM8mOBtmVJOYp36qMcULhDNEvr/b9+YsPS0XJN0RMv+dFp5+7Rj8kMP45
ltgFtZxOw8RBK01H2i0MJzLywRSux1u1hhKmxV/0FL6jgp+/ZlkhfbncZw2zN1n9lS9oIBIUCKic
/ZmoUAOO7d+3MGRou6UlJ3xU57AJ6evtk4QjU+e751tsVT+JJ2sDHyfudDrNmR825AFxv3uhIunl
Dk7Lq7upqVh5BFU3htSOOfmgqS/j5C9vGrPJKoY+kUc3dtq0LcXVgreZPW3+jQoTzyp1CGGmJAnh
63IgZjBtNQ2QvznHVbHiitbfw8WLPznQZ2c1SG/JJsZ1ytZfLA8LtS1yOjqP/gJwcARf8QR1bwB2
3Teo75hj3kyJ5bn4S3ZWzlgoCyR55SxZVShh/OmSO86DnHCZBtVQ0C6e6D7MyxtLrhLDkC5OsK89
QeEk5STILvu673ihFBQy4r5nK5PQOEA096s8va1WRAnkmXWYpGxO5qCHZ0gdoEM7RAEf17awRdfl
CeZWvnQtvtrkPCzahk3oOaCP7Vc9iOMaSVlewxMoWwzRMHr65zCa47y6+rBxrYCqxr3CD16bigyL
g2I9XrQ4DgGQdgTjjCXnWEIVMiBfmiTKISLuRbp5iVxf3H3qo4A/dA1iOGU36ygB+LnyrNDjCwA0
Z2mbMnY7h78A+TZuT4txAEMmovscdVPToUR8A1CngfqgxQXn3qDFO8ygGQKk3EnR3qB4A9OOwkwe
AOa7dG09F/4y4dfEX1Af9p7dKPQ4PrOoWT92epg5oWKvIDiQxRWYc+csrQQgEuNAORQHYgvJXDe3
qwS6ln4hXKO4sgNn/3tEFJo+YClAFBCv7Et4Nk5Zr3x8d9PJXh2vuBKyQHDe0FuuswiSpDrA9GoK
+L01t7q2Y2T+k5rBO3RLQECxCPzxDdy5R812haCgG/bccSKuuONosJIJCGbuHIbtcD+KeDmYi9bO
DmRE5uhtfM0K1pLdSXDMeL+qcCHaxPFXOhLUfeVt331V83urAUvGhT7uz7wl31nxNqGGolAmzWu4
knqJm84M5eIfFgol1eS5eHbxNoowLj7eEnGe3vKBqLmebGuSsFvHdDSgQmmGG4rU31qgM95MSGd5
ix/aT9C1B3ARphBqcxFBfnL78mHlVZo471bNRiN8mKv6rReJIx17JUq8tKXGGpG3Dx8UvU1ImVUV
9W4/PXC2n5qIyaM1WlsrJNjLOwfcETglFzSQ6nk81sgS24SdvVGl6fpQRbJoFAnwVa+cfnTsj5MO
U+FByd3smGW4yBE+baA2C04R+J81t4f6Qg27H1UA1x2VG/60m+kDaLQOxVbj2AjPjWpAMmqjkmc+
8F7uRzhWQs03faZeSIesfALd6Wns3zMFgY9s8IQbiYiszPogK6QfcQKodd9NT8X4BaqnpUM6GFee
1XGnMk9ixJWMmYT3IoqH3Ru8yBLUl9kDJJMOc9GYUMU1nbuXIvH58saYKT02tT8KAp6DLR/ifF2+
ERUYi8Ef5JqzMUJmTNM7TdMtS9zn6eFqR4xsMYmsf3O/2AAdtDhxN6cUlwfIcDqwqqTeFEOFh8zx
kKXXnn/5LoQDke6LzSYDkLxO2czjLm6vO5dq0N2JScqj1JCAMOkV+c1aR/0xlce9TXya48oaolx8
zUszOHlhYmFnRiB4MPY5cgXvFzKwuJ4TyKv1IDSDeDyGRzPts8plCPY/KcONy3pqIEuYbHxk/ZKo
SYUi43s1t7KEoiLTequr4wTGgri7Uyw7A1Als+zzyIM4D0Wj+zGhMWgVASv1qjuI5teZ79Fa1IM0
WTKAo4GiErgtn9sCI4JX7m2HlS6uPInDwtkDz3POYocMqBgPD+JUWSQo+0mrJXfL3EFhMe59f31X
iqI7VopJenLWfrM8Way0Ty5gg0uM/lVFzPtrMuBjfb/LZN802UHYHVNBksA3JTi6JiU5/JamOUv9
G/yjNgi/QbpqGAhP8VxSottiQE8CwrH5b6hkOOJSvILR0syVfbRcORwfDaXn1hcb9jJhH7rn720o
twlYwbMGfQlF6hFMVo5p/xdhc5VNoMafdBpiA4KFpXTXUyzCpu+10VbsEw1hwjNDT0FrJvob6+3U
GAUuAjmFEHMNg/d0G8dQJo55AJs8hA+Srvht6TllVIEvETZQbXW1uwyPSUxMNz3b+Mf5MNqARXla
bs0ljL48qqvyRDux1f640DjlhK9HS8VNTHkaqmSRElV5q/G8gKa9kI7hT8TdKBJtJ7fiplmrBfPl
473QlF1JVnSYP20FlK7DSCLhFXrSOxomy1O8lgUpMzAyApCPp2MhxJ8TJS8KZz8WITQRJe9SRRVS
hC5k/jfTf2KUxL45wEU41JlTMNVrURTdqNTrykPnh9WwoHOFoXA5wrazjZXSwSSTtmhdoodwc8Mv
RzZcZpzR4L3sqQLQylWoRTn8qP2iU4ST3slY7T0yukCxPv7wKVhiRkcs3fVjzTCu5hsSbagGCy1B
1FLbfqDumX58C87F0xRngQ1J8+MgMNEug49tfAh/zrRoevsDvBYGWHac2rskyoq2Qng/uazHF7Xv
4/D2y2sD21AS4HSwDOWfYIXT2SuUf40Z3yiUk/mvWecX5BERnfBHlXf0gk8VoubcfbluNeiY6d9M
v+COduKFiR1GmEmlB34k9F4qrzAvngD4AEMlnxv99X+T2ZdxVuZynFaeubGYJEhmFUpueakYfBdk
iUrzsccVOZ4vEZkbv8pY58tyZY3K+ztHbXX7LYxHYkyfpLhk8crfJ/o2gOQ5syy7WMiWZpcX1Qic
opIzz4kIeTzX41o8ROwEXDUnNGTc7rVMQySWLcf+7ErQVNs84RPXkW2kNRB0zS7JuQ+DcaQL1HEV
9ziktuefUOBZKtNL2fBSCQqGl0RfcuVYscIZBVgAPy3wPsQQ4ZfUtUFqiUcTULIU8nPZnDBnib2+
F9lqQyHkdTzHYXsgvfYDrDdvlxBts4/PGc9l+51X1z/1x8kEXwCbZRdhrnz3lCKkbnFsDOZSj4y6
JH4NUu+ydWobfyIZsLK29nGDPGYTPmSwSbGZYpPytNUG1P/+V/Ou5rBNaLzVWPiWjdQqWmFoOQip
IehZYpnWaRpJoeY5+gVTK4MAjjKrJ2TEQ+F99xM+MfrcJdd2CYetw0nyWhxqdyrPzEPaVpEOt7Dd
3BcgNzj9OknLBzoEYIAM/HH8WogoFRUDFOoRZAdJJi2urSKwX8iYuWUHYksjb5Jo2JHzlNfoxLbt
a1EsFed394O4cLkcuRn9BqcOFlJWQNO6H5BDVsXiBK/F8yIj79cn6Q1M+q2CvOGZPLfLnt7JpfXk
VBwDUulOHHXDR3QeaMWaUF/XLYH3LpsGnZlseRHEOkwWnmEOsZrOVJYJmlT4adi9N9L26FMi1B48
m5JXCYmHlOoQx+1uqZ8Z9LaINiqg+Qjw896ClJqksYWtNWvhGU98cVzSO9ulC/bSo+Eos2//RjFB
jX6OVqYOgjxkYLp455JPjOJWqVBcDInN5ZIF6VxGLCCfUdyAtZd/+8wA5VXuxH4/RU5wzY3wtsE7
KFpnGb3yImcqBRHMyTbi41iiJscdvqP3a2mWYPN9mkowiv8CVspVnnZ6fFd4CL3KIYAhS9BuERPP
d5DnChnpsVwRVMJVxrKYL+gRjKRFexQIMAE8awc+nEx7US/6Yo5k22bYKpMSxWRiP1VcA7SkpQ8W
k4LlJhWNWmQLtuUfR3x/q9fDlpA1/2rsQuuBxjLLMx7KQFza0ZW6nmZMid1EKPvDBOqb9WuXRHvS
v6uZ52LuVWaaBOVUbYi6qUg/65sbAbZAyUgz1bcoWP14W7U6bjbCmIOPXTeM0Y+EkTtQweuFJtDe
XaRlwtE5QzGW1vHknlS8k+BwkUtjAN4Lb69bHjqYn2pwvukknmR5ziXLAXQDJytKbSS0U4uIxPHp
W/t/dE/Ptl23qwROiYGK7PRms8kk20197M4yM3vNbMpAH1m22P6Aa0S8woiRIRJpwl7RqFziWavG
UkBeVFCX6rYvq9x9zf5E9KPPfkb4KpLBsCNf6IycpgYx01ZAtGLhPosEQST5JnYRnFQM9l26BDhy
Z0UAXhtC34EEvxZDeqjD6fIqcFjDQ1OBdls0Qj5H2rzSCIpRDaY7B5MngmFegCYpDuZQOw2q9K6l
44WYvhg07n0nYreeH02/+X3d/aG5Gvry2N57TIvSNngeszaFgrc+VjrkhBk2ImssGUSoEN5Clxdd
4vHEgx/lkAydL+SiPU+85P4Tb34sqIAma9ea2/bCWzXP5EAwku4ECDROXNGbfqr8pRRJ9auYD/y4
6NIidU8ptBdRzL2SA8Ewzo7iOW7jLgntoZsbci4BNOZK6RCNOtkCdK+rjAofIDRJr/r+0keqLTc7
hn/W3LoAKQM95TdKY/JH116VwJPqC03EqOwweuS5haZQfw1TjnLHNHMlyk5oooJKlKviC3hImbfa
JJZHTi2uneEUsD7pIdWhFUZFU99NZ91raxZYkWNC+iI6hA93ENk+ARuHYjEgxtOPJtjsv0MaLYfu
MksM6wg9dJNL2lEPADKj2eF6U5qUADSdwdYDyEMrYQjOCl7LnCRApIdkAnkBawW55f6rZoZJcE4G
AAeLhqzUMMEFLOZ3IRA6mou5q677e3633Evli3WtyQ4leRB0e4vBLysfwHgVThP7WhI3uTC/YiZG
BrOs/mRR3gZetkELKOjvbXw/EI5j3JJTp2r9Acm9dwEmHEhlA89Q4ls+tICOldfq1xb+VY5oMZx9
qBAPeYgLyJ2h3o5sNzptC1aDuyinCAN1egjn6zLHweBVPGI8L8wdHrNo4Pm9i7m48jn/4IvfLZia
ewwolGDow+dCSD9349jZVDnKeeS5yoGIcsHev7cOD5q7I/v4wOCzGotiHVZlrfR4UZ6oa7SMm+LR
0q8J1hrt2HLLvK+qvR5HHXmCb8yRfWD/kig6oMhkpKqQYoI2TcoOdzWb1jUurH5e6Fmt/oWyg4M2
8tAXYUPXsByOCsZKMJImciLK1A41PMB16U021FgHc+3zPvfxEQ9zzS5MlYpAM4Ifz+krpStnQFy3
fviYlXsdGihogYaKA/2WbW484elmlw9sbF17ihifOoKAObi0UhDRruqoBcCj1x9fkf+ecfPNsW14
bdwP6jbFS8SMMrw0A+fKEV9E5OJpfyLRyi7wyRgvXjdzITiBmBR37IY8ZohO0cf3fCDDHfFPykCq
a+JSu/Ts6y4kYPGCoMQRTlR8MsHUGnWqLk7c5mUhFMr9GD2rW/M/4Q9qN1d98t9kWTiPtiHFBDyK
Hqh24hzJKglvJSyhA7rJMX8CdgBLyw5c57b+ghMUQ99JmTxgKpKtRLcA3XWmIN5/wooZOg8bL7JK
QRV3NN/DTe2DmKGJjBTDCb0zJ+024Sf5FQ4T6V4gzQIMS+i2cYfyst1ONVGMQctYqTcs7yx975Zj
ACP7R4hasL9DQBDWa8m7oLRQzgN35svqaGcMhciCkFDpoXm5sfqpP9qU/lreq1CAXNezvIFVeMNo
Dw/51X9WL/bEGt3i9UCmV36vV4PtZpxoukQCmn2qjXUPMRtwyMDsQB9LD2g7PuqNlWRj3dEAG5ZB
q+eWlJeqRiPS+Lenbkt+Wvb/JCTreZEtby1cOIsWjp9VJhIp6sZ8V7GveZwsdNxNGO3g1+WRzVBa
wt5wTMAYNQzIy9toNwIbd1zt5tTx2RWGbETH4MI3qhdtlqeehuWeCupjDZB8UmM6VlrU6etp611l
kJjg6kiw/OL0AwZEE9hYriNtuIsWqc9Av0W36lSpJAebyOqWMMg+fIB/UPIUkekUCIQJZViPGHPG
WWgkEnFpcEfNiP3u34i4XJNB/yYgw6yUzWKN/eoLDQoj6u7lkz+4KtDkmCuAJOXaTuvbZ9RJGLDy
drIlBJTvWuYct3HLL5YdWccJLSUm7MDG96zFUBp2To0PGD2krCrTufgDBT0BzQ2TE+ix253WxWl/
4blwdxVfpp8g3wbBRRAoykelXxCglVLT+qt/8W7s64J4MnOrI17XP3oTN45Lfpzi80ZVtKT9mkbD
o0whqMmeBlOVSBKf2QGKxnGB2f8wDrqRoNAxlAl3d8PZYUvrtQRasbDn2V/kkNjbg/PX7ME3g+fc
hjB05Xyq7VxCcLYE5oqs9cenS5ZRwXx3UJHIO1tpNdhvMpHr28rPqFqvTC2WI0eEMsd+IeV8u5kE
vJFI7TX3wqau600ppfpXt4sbH6GNdoeKs+FdoxAArY+Uw+GOWoJm3Pp4lvxWl7Jm5U0RbktJuztO
TBGK8C0v02pQGFSnso9E5PU3Q6QbFB+zpCntkjij2uNrJ41y8e2sWIpok3eKouBhQB5KSJC/n5D7
qX2behDjCfgk6u+4Ln24SSOHcFI3LKg8WOZaBhxK/TTTPdI5TIAYvHENnbfDi7HhlRkgv4vThWa+
PSSTgjGt8AzJRt1wyFxqtxgYFXoCQzo8denoSkH00jY8GiVx1bNV8i5Fytmi71U3t5mmJUUlw2TE
BeXgTLRZVbRC2W3QtFFxSiIUMumexmctwKj04kKvLTy51wK0nBOG1uWkAj6LRIMBHhJvdWEexL2/
kND0LTUHc+nT66XGQzbrmqdtIKnCjuUPkpnrP2BAg8H7gITd2qSzPKH0R4kFjHqC0rOAUXI3slT5
2LFZcSV94RfOBV9acz/xPDRyqC8qliwHmHdMRu2Hqu2rwFPZ+uecnZ/iO58R34OQbh5ShjkjlUfh
FAKM+QM+Yqop5L/wa8aA7fRUz9jy2MJNy3e+ccRI9ZtpOUmSbCK56DgHygs6onFs8Yv/FX1vDBm+
tfawduZi/6EscU0s+PyXrOpzebSnAF6OXXJfc2L6APR1YLHefGgXl2b/mqm/oAysVP4iMCKL3QUS
JZAaC4z7ozWHRzR0/Z4w3zSOJXAQRDGwWs9dpIexWIl4Wmu3Vqq/73g95ekTqvvAssJWcZ1ffI/Y
owZu6Q8c6mSyp4w/aN1UPNs/8bPOGPy7QBQzitDoVXvuSImsjA/TXasvZrVA/N4n+MQQuaa+lbZ2
UIDj9wZN5selaAqkItkf8Nz8zJo4wi43wnJ9saPqjOhJe0Zvt6EN/KPgS5XbppIm6ATf8DG0ZvwV
JOl8lCyCFhVibulKfCi0GgOBtg+H5SK+8VMi2nnbPQPCznaqLu7D+D2rHM+yex+2LFKMLm65dGBL
7LALP7GIYkn0mtkKsRqJKUAw1Fl6bdqQr6WsC6tLmUFH15LX8KWam50abq96K/7Wjp3Sc+otKu9A
ivmkYWCJUUj0DKzForLromKYT5maa5hv7hn5nuzaC0fMjFNKXEB2Qf73Zmh8aYZg2AtNsHv0HeBl
sOoHQr8Iaepp1bFme3CNSU9Kb1Nu96WRrOg+8qbk1/jV5GC3iY0KLAGQRp5POe7cGqi5dNyLcjYC
3z0k+BkEFjEiDRsYGYT7VUyMGcSsy9+iJxrRdKxma6yQZNpApHWefwytf7IZl2m3R/tDE7SeLG3V
1uyazXhCR3mzM/J+RPU5vqupAfC9tP9t9APM2d9rdbIB49qE1AVRdddK4uUtVW9vjvPUNa1XGbwA
LRFBdN/b9g6UNiekJNuqzogvuIy4rLvGxbFjQ3F3VsXxV9KFI2h/c5N+i+saBqy4HLMEbI0bRMo1
jHXzn/OU8p0JO2K/rsB1F/oHkdQBqV+Q/EiheYcmzaAwy8PvNmVu0DbIp9VA/BCm3eoRaOeRM0dT
aCdYKnLlO3fUJ8rMVDgn/5d5TDTJpDdhVKOsTzo21/SKWWiA6nb1Y9fnxgTG1mS6cRdsw6jsY1rv
A47o0jWxLIHjv47KAr+4MQmAKZZO1n8rWWFH1blO6+WuwZRaXxvdSdvrisIGU+mqQCwimb77nBhf
SrJZy12VJNtbkQnBCmU77vo8SIB0JjtMObz5mW4TiAdMnydZLKDc37IaYv6hyGhcS0ddlRbnWj/N
Wafw+euul+ltiBZlnnn1pPZj91rkiAqrm/O+TO77k3Izl81NZ94Fq1dSHSywhb/bwKP0RvmC6c7e
APfoCIAH0ZFwDjzc5YFLgDOkp5mODfazwvLfAde5cVghtpXS6kicjQaQ31RFI/61mjzrI0fqq9Pe
i7K5gy89vsFSfKpbHNIpDmOqm17K3gOTxWUOFlmudV+/0QiC8VvbKu8k4ZjczSMCvOmr3Nb5c441
AZte9Mc90KwxW51bWPteYAhOEQmSi+HAQB1RuaKUMVvK9Lw9FEN1ykw82CofKlFMp3eugsc88Ckd
hx0Pa/Mz+f3RaQLyImcXU1RIMShCU/Y/hJvY4bkzMYB9ZsngXioigy8Z7WHYGXOvYJDbZfeP/V89
0Kntgj+lu4Oa3PYtDvESCk7rbMysaD/itaAAR7NjFA5LtpCeO++l5PRAcvhYwbqK16CpwHqpgQ+e
P2nQkdmo78yl2nuSSIgTSjBED0y/26BzaTSsHzc42CcqedtbRLNtch9f98SBa86rPJqzHMR1Gem7
Nx1oxG+Qc6Mt/v11umds67ZfsoPqETd/DiFm+y+brvR1njT6AOr4lESNZQwyXDVc0NTYHxCK2hkT
Ez+55JXhksaX1HqyOYXvtO3dUnQUit0JJfPWMEovq64qBS5tC/FTJGuxEVEJSRrnpB4ZCCxSJxED
d2sAnln+vZUhi0TadPAy8+s2K+5UP5BAxnMCi5HGjHD+IVx7cI19DpWcOXM+EkY6s/dUHbT1iWSz
+440PlSCchtfGqVxT3V8k7mwQXpY+2dBIQhL7BvsOQtL8FTlmcEiyZxRPii7JOeGNtDa2apugtDq
9AnzNVlaTFF5yiBw1bgcUOUjwXGzCyp6QW5mUmxNro2jTY/cgRNhbE2LUzcR+7GqtOIDsrdIScOD
y//MYt0a8NE2QDev/7zsavbvRvPRoe3XjgasQ0sbogbctzdrOAz4krTWqzQWM/kGmtt9+sx7PLdw
PbSyqQqmp9qDvneEmPxQkH2k1q8hedJepr2p7nH00pg8w1fcOmhuQI6IMCJQqdJRorEJ/DHPCjEq
3s3n33ecdd1nKhkE3pl2wXOlMn/INEwRcDBLilki2dQxlj4jZyhRBK6ya7y2uM0rsEAd/rjFRRp7
NstGjhO1CkXVxaOI15ox3M1/AjKpiV2PPxhUK7a8Z7k0/Bj76xp69TWyas6CdROrWl4h7bFyPb2E
FN/Ty8ABiXaHaCr7AtG3N9YbxBeFlT36XS/bRFISEvnVYP7sQwBSUsDXx8C5CmCyx+LaqrSQ/CVy
SbGUeXCL0r3fcaHU8b9QhKVPpjcATuCCG6w39djbiYKaC1kXoXjsG9xVt2KxKE9q2ie4aswDPRQG
HAileTlKzkXo01w5+MTVwcbEVc81ImtAWhyCSnWha4zJ0Rfnu0yv3WS7zln5Dka7vTvr3pwa1FH5
JNT8Gc0J97+LBUt02+DKIlXMPU0N1zotSr7k4ljbkrNq2Cn37xbbAEA0w0McaY8UybilkLn/jjf0
klmdPezW1HCVMbKE2EkvKF1xsy2JPsMgLoIGK77z4F6uXt4xpORIyXQSu/5irlLakW3wbMwovKVP
ii8dSnrPcLmG0F9/z8vj9lfl5Dyo7YBS8zBv3a5Ubd+2kE252fdM40ugXN+LkromYINeHvDUgv7g
VPq1QrZDRB1DlJglVKjItvcnedzgy624UBkQgKybz1wXg7xbMQ/WZu4ncWkiqdOQrxQSqkFVmftU
2C5FSif2tdyYp9xUo0yuCdM14qdQ80tMJ8UbxHJDSnuiYhuotxjrFePKZBUtyNmfvWkTYPOX8VTI
rrPj4EIm82PEMmqK0AO8BbNRnBM2x+YFmSBh2+O+oDaAFtwDHlcpZgnNHMkCw+qVw2vVLPrmByZI
AR3q2dHiBdrA5R/8Z5EMIwi9kxnZZheBXS9w87CBxPUJdUPYFEd95sKb6GmpeNI5z3nFnT5pcP4k
+q18ABi6IqjUJWzhU8C65FyEAmtorkJmA9GITTwtUodiuBTHQLKawj5lglyxnhwPytTeD9Xm5ET2
jMO0i+zeR7AA/rwGdyM/uR8jAXsuSP2EK5OKCbJzNUQfZalbLDLiEsh5AP7k4EL1Ap8ai5BB/N6P
98R4Z37al3Af3DPAarsrUE8GKaMqYGokwx0xPCWLB18qleelpS6gtObfAnVz3DdM9WWUN8iH01hl
/WaA+D6qU124l6Z+aRZJ4EDD3uZSqxhMsVzxwmqsejwDLh/vIOc0Nhz6wJioJ36rROG1edggYAt0
+o2LjJf6hPyW7xcKpnSiuJXFfzLbpA1MveCBQjyvX72pIhR+zJqYdo8mUPEdvWx4bkDgWQAqrs8u
Ya66XCmXw4dousaSwm1+9W1/L9VbDZsvioqBGYSFSALTAe89JtmIGsru4NUQ/FIjyeLH9c92XZQj
1mUj8ErW2eTOnMBMYz/kKewJDn+fCfOQrn0Ff+9j8MJcZOR8ab+wkzTLTvPo6zgo2zJKbW1Bl/Li
+P+WxgzBL2XgwXEplsDXknVU/ANEjiWa5IlYi2yQ1VnAZVP+5qWpdTTA+i5n8jsxfmk0HtfTPGQf
JKaitam/QEOLJRj0fwNps3I3Bht69L9yxKhdf38R8nIUDWwrOk6SLy65nECcoVxl4EfFyJWwTdP2
3NeVYY2nZuWR/aarcESLLkqqmnaxdckcdHqsSj6QS7F+pA324yXACRb+wwRek0DEZvA6HAj0RGNN
4cMR6uL0rfJhvRsMZV7MG51ZIwzAIxtLS9vZcuGti2tJUgAAihtDhVGBlP2cXh+hFSr2do/46RuT
BxXs3R91gdTVUvt62WZIuBrz5Q8eF9zxTTbwEAzMR7Wk8MudJaCr/0d8A+bdozOvKktVWkIIjfSk
TE2b0QGQ16EM46x+EicXP+VVGFYY/GNO0Q1iXsbM3UdF6jYJ5ss/aDQ+abz3XVR+zoaErAHZ8cdA
VE1ua5RPb+m2kdXNuuQ+wafjSOv26Bm/1jgyoQ0miCqeKhL6kSv+MKmY4FA8xfC82xocb/R2Lwni
nWltIhQmBOmgBDAkQ8q3P642Tw4neo316UacLYiqGNH1m6iA3D73hhbd9bteJe8p8uVntbcgeEEX
o+L1fb07TfvVMaCHc5FxorjIOGFPjoJFrHFFqfV/JeQKl14m1ScZxpWnTeekhFXvlNqrkAP1RF3o
qJ+xhQM68VvLhoaw2xzLleR2lCRR1NMVNRuldnWEv2VAYz1hdmmGZ9o5Qzg4pfFJ40HQ+6fdQaEY
O6bUAnVgadA7cYQCEiLiAyTsJ3nOU9Kmn2XLz6lH9PcwF1fzR+pJp8gd2neXaVQ4xucOpl/0Z9L3
zDPUoi2voKGhb6GFcvEOO40Pyy83hYsCz5Vv6rhgy0O21Bo4z258or6Pky328m4eXPWU7W8dKH1y
WrWleet0KzWZqaIGzKTaPf/bqCe79sS2YadxPFN9qI6dpkkovMAQKRm+NmrvpUVv+079FuGpqVu+
yF3b3MtFUj+jFclfGb4ZjAScJmipcv26g8gNfg/NcafZ5575qHkQTXnKb4f4EX4Nq898r6PVcqG0
JlX9rGpwxKPw9wHlzcultQU27nwdY/ggpgddTS9TztbNnou7jtAQskR7LiNxq1wFhFN7XMpqEasx
ZjHBNWQseD49vXdxtrymz2JmoxIf/WhUVldV/656aJSLaSORDFMh6/FB2ZBaEwhku/z0PsJw5sbU
MQv66Bfm85wLvCLnRYdI8kSDdBo8nNxt6glno+1YeVQJ+2U7Iq0NzBv5RRDD6YrC9RoNdxfjDjy1
+tQUOLLFKnJfvUt5snWVC/aElr/5oT3gooXTuuC/t8VDBz/Gkoc7YgKadgT7DgdgGyfixGiM/I2K
Z6Xe+oy9rVIOAeTHG3H9TFx6LY+F/As/rEDLi6cS0oQ+udVgo997x2hfAzX96gGS+XXcC3JxxqIy
ud+XijPVYfJbaBSrBNezByfx60V0ikmygY6cEAC+QKdpe9b3df25MomSGmh4AGbw0oxiv04AjNkt
QC/wZ/fJnuMN4+MMA9XFimHELNVhPmbBOv08ZvznQB7+qfOq07yyfLBmW+7q2if/c7lg1nglBGFe
z7RZ3RvQda6K5JewXzpZCGHO5oOynI50aENPRX/Cjv7fva4+yAyHNqV+GArtRlsNrtKe2NUHZOa6
mdqL2ugFx5v6sB3CfewPj03ey1cNt3YiE6eQ7fv9XVaO/mGl4Jb0PXtb2WyoHVPBLz9a80qspPe9
fHpB6ZPk6PQFxKuKRrjwXoHnrOEhEiWyUX9gQpIWxCFqbVh6E6D9CW7P4Q81DnPJuXxtxSmtAH7K
C5gfWSTFHDmDllLQ1k5Ry4Tuy6Jsfw0L6KTeUwkvdqRCThO+jMO10lGeXZaZDNNLB23VxZE4zzc3
8mQ5e4KtdU+rTFxCzrSsHbxDy7tbepTuPngq/DutXtR+oQOIurB+RGsvtAP6lh7bmM9wlXCT3QzP
j+/LzsUobRVtgpULxa9oo6ilckGvAqaHpsYJCPzHjSU9skvsZ8SC0DESr3jHEhZwxa4oYDEk3gtG
I2gnhbiervpwjTl8mYGQMQLL+OMrEz1UNWG2x45Lek+9twmmcYmC34G2Aw0nXlw7mdJ7js6DCcQY
VzQV3SgspKObVqX2KJdah6RIhoJLid5mGIEmPV3HRCDwbk5MLNMA4L0LlYBLvWpaYLy5zmn6de+l
lvSXTndbJu4GYjsVvb8oGHS4Exm+OwFOZrnCBc+mM9Tu9wzgNd75IMx3w+BAmMGm667PapIzN2kB
7OST8YTocboFEl3T9zVhIbZWdjpD1wYHsM97/c8A2LInWRZSCIKtCH8QwQ3W+Mx2rSXxQHRYSH9q
82hAv+GVL3MRLfXbrfYF2o5NomA8XilScsto/7pdJtSiV/YdWdKkWC53VsxoldU+RVKH5wbO5nMY
QxignaaRjq3CnSaDgBGZguSnMSZJsPYT/YP1DuHDwt7IOCFqo3Kf6x6II82LTNd0AFOnvamJXjFl
M1zb+eBlpuW8Mrv6j7i4t3lkDIEjiCbRmCxFJXwM/G3pB8em6IisRsB85nUmfL5OoRaL+DvXIiZK
Cng+tNKJhxA0cemHAwkEPk7kKZjiX9Srd5BLu9vlvUXlMKIQqnz8glgS2BeYw5+lgLdML6aEAJQC
JZyEsCWk0qV0FRRaly0Ax7KGDNeoL5rukLXtlnmPlqGIADJ68J50jd+pLEi6xa+Js1meAbr7d1UM
l+RxNBbm+vkIIbSF6u3zYJSW62thxwCVRnUxUmWio5KxMKKwN+grriqW/q8PzsaF9G4Wr/tVqGY6
afcf7CvbQLBjvbS7KoM3O9q9r3DSC40ZlTEDX1yvEhmHHLYidXuK9n4DmzqQ/rc1nd/VYmcZFDA2
qzFm4Sr4YqoEn/8ZOo3PHmu4NqGAQfnZN++AQ723pEdwdU3b2lDpDGGlWe10el2p3MPEIGvXv2Nr
yZGuahJaS69h4eEi8JTP5iLZ1GwniNKX35tdulpmgwlzTQ6p1iL0IY7YZ+aer0RBGybannd2Lqvv
/Uv/kdz0YK8O8xmRTCVl988FKT10n+j21J2hwloG3nSyWoZPTgp3QAXLqAHwsA8BealC+RAwIAqs
wuMYU6Ys5WsZYIzcxIbwf5z69TemtttD7nUuCHKNy0B5FqP2szsEMgoGwpbUP0Xa0gSFLB1ufq9q
8JuRQYXZkCJaRWWwxsP6OVUk/wUSyjstTM/lQPIa0C1c+1cza2i8k0AH4G4WwcGlkXNdZd2V/TGf
zSBBzBIfYGXHzi/Vp5987ShOhUGRVxRlWHU13DEBtRAp58vDk5Tav4jNIJG+DIrpZeD/Kqz0URDZ
ItASosF0WoB4Ilv2y0XZLdKwu+1TTbm22XFqLSD9tTuebYSz3hN0wIcxddkBGOkn/34Tth0GUI4B
nf12mpn/uyTMPynAPvegzCsw2pk5mQqdpCjJlV3PP+zT8Ys4B2ZJAGuORtlZmYwMRit3Iq6Wto5W
ZeGjmhPszBsiQCZlGvPYjy+5Gw28sGkz3KrHCbGfwddgjmDGiSNZw8wF0lV2i6KkKGBSHhZapEUh
o8ua5rqy057DL177cnYt8sBPE31LJcdR7gmqvz7N9lxDHtNPDYrLx3GqmJruKPdLmGSx374F4saP
H9Wbz4geqyxipKRU2P1xvz5Ma3dGp5lVePPk41pBb+l5PxEWvX7eNLKfPX7zsUPIE28w5/TXxF3x
FgxOn7euuO/eUWT7ZC3lkb9WtkArbGcpO2cFRVu+GTMUP90R433LVnDJIXvov2V1SSSVGf+3BOvs
V7ZZbhFq5fUUAF5M2mNteyr+3zDfQvJZcPhxGx0703dTQIC8lK8b+Ng3yRIOZu2XiFDFk/y+805w
UEwmsVKysD7tVbkmkPI/CF/SvyJzT7k8pAeqkdpncydpFvS3gBgB6akmvke7YLy311L/EB/9Xlrn
5Zu2InVYNe0E+T/pU6X7O24dzmPl2Csgb/9aGVHpzZCI8CofhxmEFXTwgeIN9+XsFypdYKk8FedB
7jK0ROIfzQNrgtp+DzITOXY6exBUzKbI2/XTsrXZcQ4bCkp2AZ+G10LtXZ6kLcxNTY9kOQonOkIY
xCrX4PCIRdXKQMqn10Zi8nx6yd9Gm7JItccXZNRCLoSyad3ORytZDgEJojElDnbgvGXWnrBDLPQ0
fAxln7AOhsTRBUMRrqK2ya9G6AnOvno4pYB7Gd3e0X0f/+EJLnt3SI6K0mpDObupZo3rpxtrYcNh
FwwokeIkXHN0LpMhhmY7HcfHA5ujHPjGQFwn56jL+7x6jFrkIA2EdKRdXF6lXuzhAeGIpB8ukuCK
6/XCu3jY2PJLmuQJtfZ+T4gvkcCZZTDUaBsK4tgJpc8yfdSVhMEN91S8alhjYPlZHWxnYkhOZthk
bIxVjCzblI0ODQPD8Pmtc4Wl6vLjA3fWMwjmtFbXwHPHJ2mza5gXTV79a0EViVDd9nI/Nuvu+CSY
+0pe+rbHo1q+r6ee1tQ3R9X1gjLHpG5dEi2rJDDE3QrQVWlqffO4vJseHMAtfkP9wWsO8qQqGTom
BSFmRwnw10frtSoZm5TggaLPI1QiNUzcdmH4fuDbZkX8r4B3vuKXIjhvVbtiWbr6P3hPL8ssOrnS
0HhG7SDt9YSjVibdTz6XIt2DiLfRpdCIUYXsdD/q7QN6xEE3I7AuAA5W2vi2oHLkn6MlucyAZoeZ
4DqAzow1KvgSds6i05QR7m6KAAIv0vV9hdfZJEiZnlYiAaAM6TiqNyVqFyVWDUi5jA/x/nIpA1Ak
/ctdBBihb2qTJ+aFamtnVu+TYawA6+304xYnKB5kqDVG/0+byrzme80bxHXy9OZKXgJ5owdSUjaZ
xKKB8d9WEKhmoqm7ok7xmZpQQF4gi8aUO/Wt//MeAY05j4omolWL2Gy5xL+sP+2L2U6+wA/CSdqc
yS71J3Zi5kJiIuujkpMDGdsjxhrz/V5Csy2G0klceDSlScCjaWrP/vohxqTyQ+JiCYSepWJ3v87f
IMTADlI31TrrlfFHfjgfa3RGdo3mgSke1Fu6SdDUaOHSMWzawNinrBsNc78MDAq2Hr1mcxXZ1aiP
BpB2TYs1e+KvONyp2IsvvPlG7PgKx1hAMlpXOAF+aCYGa7eRFJ0QuilTWV/mikML648KJWF7T0EI
WCcflg6QNpMNLx1FXEGqU54nClo7AeB5YpXVTJwnwI/2g2VEPtssyzPkGXB34sQbD66HXVOPTLza
zJpr9sS4PvdqKMpb8cXv5KUvjL+M7W7y49BXxXAzVGGQrcYTf4qbjcMFnt2eesfaBN51EbhQPwuy
8gLQTRf59Z0phBp66Nqx7rhA7GBSxt4M6ASBWCuVacvHlEMmxgR6HaItSJ6rjhHx5nlEecC3Zjx2
N7GzreitWFhVrPqRXFvVP2vMbbV4pIVZ4QSrQKVWIdxriF/i+9tD4Jhej8QTB1amZWkTBGmOa1+d
15ykYoQ4vDmJb4g1hqBhvnWYTKasthFOa7RsrjATIIzMFUEYwMqmsjyulmXr3VYAdxnpsQzqc16j
adM88NVs+6r3dR0uX5F/KqXy5PFNzVU9v53Om4/O+OAqmGbTwPavMLCLJHSIhcxWQC+s8WpELqja
mLTllaex9qKVIhpAy1VRvrU4HXxw3F3KgY/JMRK5MLDhkPFef9SmMftCpNsWCnKCBOlGG+wAkf97
0Q1a+BNbk/sR5+mE6OkU+He2ufqitcwzT0bzRDL4zNbRCskBjpzLdv4rz5Bjui1OF2sBocEu/gQJ
zsBhkou9KXdTFdIcxsTFRoWjkGwoAm0O5b/GWolmsOmxP8I/Iv0h8kn0l2S/w0ZMZXDQfwOfZ1jG
/rdiKi5iBpo/4yaAPhGZlKUepUWXkKx0VWD5pSuZeJ22HTyI9YJVPP2SpQ+W/25o47l1kxbCzRyL
rxofjxnf0dsacj8kLxi5O617Hn6v6YkJdGstS8ESTklvVv0AOx+8lNGDP8T35hQhuGjL+ym4FPkt
WAV+tzwZBq9lmWYe2qiOR/amLU8rbsWXsMiN+zu8p/6FjfQpMtyzxXxPvLEgBZHPfVE4hSx0idaX
2Sbht9dxvEUZxL+opEyjgC0jGqx1rXFqMspesu9VXnG/2WDoxduQdlR0cukX2RhEhDcmhZx2aNIL
UwWgRvf5vOJJWBkeSCXxE205Nju9QQ0bC6s/CuuLu7yoLP41KzbMYIXh4eoIO7d3r4Bky7XFR9HN
D2MAkQpiyF4Tw6RPCBfd5abb9IXNyQJ/4sKeIRaQZfngSmAiX6vkYizepg7sjUmh9JVi86788bTe
Ij4ms0djBYINyddpIl41F62CTQoKjD0lZBDp+4WP6jZaPurP6EYGaOtwG8t9rN0f1/5fk93OBRBs
0xRncxDQxjslVGzRZvtCjYhqyzVeGFrXz4zfW0m+oTpHt4iSZHKS7aArT/Q35FGz61G3v2snKNyU
MMO2y0WgygLPqH1yENRHKLif0dlQ4YeJ4oXN7grFkTNyRxJqrsKrJZrrKp0937gHEC4HgGxSS/Lp
FxvhWlhFc5aiQ/OZaoEvBWgt+Y2Knim6v8FKD5nKzTvqTORv5xteda0ApcLaViedzlVLiye5KFg8
GGCzDDi5IOxc+cttqYZnXoctgRFI7zUFxC4wbggcM49pkUIL6TRoSCEOJWxZGtxaJ73mqaGPIX4o
MAmgOdmshAgZKpGkcOY2VlhXbibVrudczlY465XMK/13g4qnuf5mH5n6TVJmIAdK/mMud8F+ojxP
XaMMTvq5OywyJrCxZLRKxUKi9rE+crTmtPQlc5qbuiAXT4g9tdd3jt+HYfJzy5vrVq8I/Gj+7yYQ
04g5fGiHVcpMsfU/38wpu9LbEoTGiONDbSQ/qgBsRGgRVX1su/qy4cvxbfVmrWDj8GQh+ZLdMy0u
IZDFttDdM6sVFX6RPgZ7JtV+XM8zJ9hZhd2QrCemVzw80xl7zE36tvVTzBHm207aZ8wqK2ruBOwC
nv78TxhnZYuHe7CeH9BNAQ0wpVj8Lae12HDQ+BKqlFfQR1OY2b5vN5f8TVmPXGLEQA7e4CXbhHS0
Y7DwMmpNuSRG/zm2YA/e0o86yVyc/e6hkczWUmy88gsuxTEb+VV8Au/AGYzibX4gevF96bZsjJ5u
2JQc0YwLqS5d0gyZbWjNUi2Rc3qas4FcqIXOBrpiDpH2nlwoH+90QhYKQr4dhW/A4P3GbH45y3p2
ptKIiOf31RQCBIPDpOFq5Z05rr7eO6a8Q/yD9TCEelkd56QHPP1CiXC2KzdwTte1I2hhHIphMIUr
iNsAsxE34IrlTprdX2JDRL2qh6V5iRNB3rTCvgJysZHNN8H2fhNv2u1E3jTeN4coqb8SM7rO4V4D
5/mBKUIe3jf7pVjA/dc5MQWPPzmXO07u2ZAMALka8RDU2TQGwNDft4Q570TmMlTIre9Ii+0QF+GX
qDQxysuDoXhZfNQkPYIVAxt5TSSJTHhXane6lhFVKYYJIWRO3OjvSdP5eKtvJH/h+g/8+nSuEFD2
lRqKbQDaRJ0/7AjvyGy/4KCIDKGzEHnHj9BSmQuWs2yM9MDV6PsmhTpnnKsunzfeKgQKqwW6+YWV
t7NPw9JnGXGTUjTxwlVpX+TgeVlvg9M/g2ZyewZQPRh/OjDpFwvhMGTGvoXZAS1psfIa4GfX/TdH
g7/xdiM47IRwx1nC4fPHz0s6y3zd5vX95taMQ2jtllu2MutcTH7QmvbZoAMxOcGXg9n8a4Mc285w
3AI3c+l1EKj3jP019puq1plf6RfKCm0V1NWmhpUvAeOO0HjYiS+YoZFb0mf8czWIR05Nr55IyQiO
96VMAW5eRD0o1BJej7EilLyifR2HWNHor64tx8Fsicjl2aco3Q6GESn4GSSD8CL9ckBaXkpKC2Zk
YSv6AH2w4PTzJX06ZdE+G9vXjBFKUx4BCn1OcLTtNJA5MGTres/JsnBtlYm2VVi26CIXh98tQdvc
Gz2RZjAx9sdeujmAbD4ejK+omefg7zV8iPCPJIc0crVdwSykS2T+lunsIEzD/iHEhY20NQsR2GT5
85ytkPoZH4w0nWMCbRcheuV3/cIaL4nQG4/L7eubRag5/E713rlinQzbweIlKKdxG+XAwexl4q9v
Elsz6Jl4Sse8StbFmX1kWWd3BfSK67LMex6te2TSoC1B4/1+Tpy/boSHb0bHjdthWhRjo2t9N9tv
ZmUG+u7OHgss2S3zQlc/N8ml2LNs9bg/GkH5V7Y3Fz57r4zLqeCxvEArMjJMVNI6MlrPEjz4N3lT
abawkRazq2qx0d4Jxv2b2+WRn187Ig7pfHSL/FXh1c+pGAkZ/I26EkYNoUM9IjrS4iLHkRJ0XPHI
NZoJKJoYeGZn1KEWD27P9gGfEyRSGqX8YY5dQm7MhFQzec8IBFqS9RxGbfkfKP17SMJ5BGiYyaEJ
GawZiUHieJi2GBAxe8T2O/D4LATbASUmUqT80acuhyWgWbZSfVQ4DGOK1HrTxNuXK5g0pqZtN15j
krcYw4BtGcLr0OOmKB576gUfTmsmIXZi25BV718SL1SXIBUduDjGznX4B5T6vKSQF20fAaxhKw+6
WYo0RspIF22AjZi5DwpVh9ssO5/q5B5DyBZo6ZuZPXAPXe/0VyMvBrbhqOjZNhdPlxyJ7YJeEgwV
6yyLVZs40jM9I+YlFeBFxtWFT1WkldkMgc8j96FNP+xyXYWCCzkEkvyaRTRt9vxslTvYAJzqpF66
lY8ax9muL1fHlhT2/8R9zrSFL8649xOmex8KsBg+mDh8U3ZjHIF+yvvt8xvwqAMmcbuib3fvb+1s
IA/EoroD/lKiR/HsFi7+WiLREztAmUtd9vSl5hnlMAanT3WCEbX+XV3rfKANp7DNskYWcEQZr2Bp
IzmyOoXmG/dWss0cYaxZDqNrlOB/quDNCKVZmOZijX0SxjfHXaszhdLkHmcr17oxMW6He9yb5OHH
XeyrI17wtQyX+l9MteJJLt5o1WqJoCCMLIqhwze87wCtAlcCoyC4YSFcqlM2MlgnmBZKUrmt9y6h
7ji9NFwtDJGzc98RKIyha2Zbl3KJY1srUJf7VLTv9pV6usxUtCLCCf2AqWri3ZyU58tXYlU677p4
I25UnBUtrmz3enVqIv/SIY7TXU56HJIpL8iM5HIiqFkEisbtaOcCfofM+IkW8qirhiCGPDu3mxB1
gE5vuU7dNe88ob7M+PBwMJ+KldxZ+4X/Gxj1FU5xmsQPbxBtZD2A/DIF8aALx/i2VXy+Y1P3/MDc
SR+iefSDOxNNvgTSBUfZVpn/g9peaRQRdvRiXoOYyYaCRBADiYIMwnYFkvP/MwWWytWZ4mcLycVk
cO7QClQ0FMvLcFJvHhqdznYygoJEjtpeTeLGdTUt+cn2nitd2RZYahABE+NpGhupP4piaymg863+
7UTxP78o3HIGexSYFAZOezJ82h1B03GBAI+LnQIvTMV+XFhn8JoVpuq3y61+IzC5hhnsZ+ppcJxq
ugI2+p0dyZIV1hLl33+6Um3hUcxHj9bjdpqUosj5tY8+kDEVb3kuO912yr3SHWZiCU6gM9l8WTKq
2yettuuCBEYU841xkKus0TPOtTzqPpJkBQ1zO4rJ2S0y8k7lgIgSJXj5DM59G4TMsUBftJ+C9N4G
uzjFYXSyXkbDzc4NGRo2/uyrwyZajhPs7gBjJISmRBW79fGkwHpIbRFkW2vbver1TJjkacP1+pES
nCgzzhc7n+1LK4v/WRqWWfJ279F9J2RYedmW3Qm9dqvy/zuZhPCaUYSZKovxq+JgcbLrY/oQAsnI
BFleuLFfC9sjfY277KILFhiTga2hUn8swFwwi+USTGQIR+fYBcxFaCUh7q/4fcwvGJZ+/nDdtJ5R
DXhG4zWK88AHqWqa1nlXYtrOnXx1Z3/xMGOR6tyKKj+fnFkkDAVFj1/WL2rHYtcuUHWObCaN2spR
ixb5PWdix6k0DOzSdDc55v7ByBbFzvN7CJwJiMdAi+B1iAj37owcTHb3uwGzqhcd3OHHuB/I7HgH
Ef8h/H42cAxvflLV81LFI4eThwg7k7dCnfOP/Lo3uRl1486dYCzqp6tVy98ho27wPMboBttQuLi7
c75e8e1WJmaxz6moObL/ElS/iLXp02LUpraSCXkBbhOlwae15yUIs+q0pJVO0r5X8HdjHD71FfLA
iY15GvDfw+Sd0rjkF15xUgjk+wPWCPAFJoa7N2ECvhy1OgANNIvteX7hHNJ8MEwO7KXvwq3fRUw1
Aq5F8h7bl9kTZ/SDVyBWnvZX32Rpdkr6yQTtfDqJA+5nyq5kD94aetSutEFAd8e+vnCB6jWSBl9L
Yl3cF+GDENf36ebyHAkUNicX3rtkFp9G09DYmuf/8+zCWP00hvQHdDvReppWFC8Tj0+3drrOeMGT
zH1SdfA32xlvHPIgfGoo7Nh5GOKyOapHFaE60HrJbm1qTJyAPJ1wKWC60+V4EXaBn+wmnUU28jMg
93pbmhF1oBvU9AXDdi3xQIFak2SibgWDk0nXNHye7OGp2wUqoD+0DeskZ6CD2aPsWVxH4QblRis7
JTH0NXoeYYy+Yl69HWxoKqk9wgFwEK0HTlPo+N7zLoP+kzyYKpi4w9YLyumb2TPvHVE3nw3FeL2k
oBucX7vJr9Dbkn90iWHV02x+a5r37saQubIgIhbW2/Ic8iCaIwx6YZsl2yeEc0cBVyXWQal9CtU5
remv6ePyFoVc0Xjx48XOdhYoA1OjxnaEVRBWDCHvJ4V4CNnTBcALfL+Xzo81xbZvGJ306LmGYBsl
MYjTqpXVDmVDN/4tRu2CDviWCvWgjcFDBS2aFOJ2nA5HCR8ilcDjtBcTuL4b9wnfgPg0miVpdGlf
KKKQx6oA/uDPde21+Wu2m8d6Ywwx1Ze9am9b0C+unQZzWdjttF5XgDKRW7WQc42iQ+4jt8MDrqNI
5WM/X4C5YBGN/kCYVCLTp6Biq/X2x6Gbp4i3h6h7SwhrEwvJFWS5NdZXip8P1UOAlWvXlUcfzNS5
rgnQHr/DVuPxLGSnSn6ToTJLI8dCTf69DIb6+Q3fTKQOdysEc3nME1fx7QujpZUrCGuK/9iEwpy/
ZEiAAs8mOcsruwI1ZvhmHt9FfhZpe4uDhH55oE9cT234DMaNQhrsNTjSwtf3zgzi8VkxaAc2OUZc
Hj3nNosmZUpYbEC6/hgYkfML37Hu8L5IWNDQrc4YMqn0cfYW1SasdGDAOyYzIchFbJiOE5/GuBY9
tbeNBDbl/YI9qj+7MowS5KB0sg7iFOueCALT310ltWaLXfAt0xdRQNNVe7scFvPG6Pf1mSTBHZM/
QSEjjlxCi8uniIYIoatZZkPcqD08m2pMPJODLhb8uZkbYsDtwgSQy6gLiOKVyEPQVDR/ABfltlJL
ZpD4wxAUyRgnius9iE2vVqhe5FCv4Gr2IRJOHh0U58alp8I/7k+4ZVVGklb4xlKvvT1goLg5rt9H
C8dmFF6WxLna+FbQ4onVYXdPaM2FH92pCRYloX9+eTV0qfNirXwiaJqqtNFmmHKBkP7esbkjxbZ0
E/6xH85espNANW6bhyqCAIykPjOTtNMJ2KZbMgPZwE7gF+dcPePN54ckr4dHQyY3srAJcYdyvjI8
EkzdiBRhfEffxZeYWBUmzsRQTmafT9IhDxY7meXsEdMCrO2XW4KcVtEYwmj5U4a1RHblmSvS4Kdk
L3AaXfm58UzGPAoVlcu8qcGWetUGBxwOYhIT9dle9AIgOWWnpmVFI4OH0F7YJOkJ4Yq3ScZDa3n/
PaNY9yyKTnEQ88reaEl5TJNRvZlQdg+vQ7DE1v8ASX295V8S1JCKgT6yKZQp3Q/EQOeYMwBD+YVX
A1ksFAsfWopOvXvhiTlAGl3RCZP1jX/ZFcX8CWFbiz1HZGxvgRFSovx52Pj9fdXDY7/fT2tF4499
xypN7Ys6GqTZxszIV/Cr4scHKtCK+pLPToWoIgvnBEKCWBsESO7nvSafwFmraBBt+vNCaoYMKGlZ
fb26UtXdstROZYg7s9gdEi9WeLd+G82g27T7oqA24/yUHqWvfu8QbtUCH6D0S7Bhx/olpBRoFS14
CELTuuEWNr5WGR6gevC9SrbkR7UUdAWfvVFR1Iyh/JWvTtHBxsCl+mZW/evDFi6TyZ13bp/Fuqvo
Vmazs6KDRUzUicGc/utBfBRf2cpvAQRXYs9zRugKQhz+5M495Mk6pwwPX2r4I6v9ALgVb+KuzlPF
2MG2z4FcUBbvJmTD2dtOiuVFcLfYqOTLRrWrdeRud4nIy2JEJGGy6eCityWceH5gcN8JIcC7tUR2
7KCWU9uI2pbz6/NV/he00pzUTKszvg0JrgRZKICIL5v5L1Rs8yzs44T6U7a9O8JUftZCHTugqdau
3wHvoQFPyls1DdeGFw3oQeW5QgQ+T+rf2NZsatwTZilkTp21lYJGjquG8Iz0jNmNfGYDmg+maeVl
ktVJpkxgrJU/vTAwfMyFK5BtO2eADobFn3z6cR/rbrrxIkbC40mBiNwDOaBU/UdVdunXahMtO4ov
1r9R5C8qs1UgZkqxqzWFux+s7qoWsZJ5fq99hvDummgvvYupN9a11Mm9GfgqFDEufTQXVWHNoF7i
xKWGltnaEmgpTHOr9apO00uKQuF5eQku4RnCrYCuvRDEEqglIDV/hYiAZ1oTSnsq8R2Qc0OT77/C
7Y9PDVJUseB1o4P7Gt0+LPwTkwlNBCoJ1YO6GXzKTLhg3UpsStnt9shWbBlph+0X0B2cwA/MSKKl
y+aOESGL0p/CHar5k+FdRzY0sdH3KOjfsjoqSm7va3weZiBMIBFDZaAWyQE4hRYoU+wQlu0FJrWJ
wTuDE4pTmjzTLaOkgMdSr3lfS6Z4KrEO8R4aLFHKCCzc9B8AD+MJiywtSWAvPatmvH5wR5c0lmBl
0f62Z1gGOaDMU+RCRkEYlzqiStE2lYHtlcBy+ORhfenBrMJCO1Y3JjS7qfTk3MtT1cZhhHR1yfVa
dDfm/wCausjzsgQoc3cyvHhXlmE6bSxol9qkrHNon14LgOsrdabNjryUnUfT7D8y7KuBzzNIw217
7/MdORRjdUGsBhB5WzN4mUXqZ9SpPjrxdLRfn3jWXwCCspf2B7yRGWCGeb5IRnp8pmrIU5RIGW5C
hS7mBB7dmsNbS6qLzo9lRu42nfgQezS27DISaCGkBuve/TZk8AoqY/2dr4IQCaGUB8hmVKbPPZz6
VFvojn7cz03pbOPRkcNNO9Chbplk/sc6wp+AJN+we2yCeU6sohr8u/b2FGYO+oUoj0XbOrSD9PMn
8cpxpv+U+LbBgvYJr8QfbUMk7LSmQsBByDfaBc5anoqfGrg5bz4T5eQmX2CZoZmn8z+fWqOFfiiK
zva/U4PFwY7NEo72YCtM4OEIQJRK2J/TWmrSMG83AY3zoMGgENv+DtApy9B48Ts23wtPOAfnmwmd
stoSg5/uY+8JXZOsTAD8SVhbGlkRgkHauyTKxrvELd/pBeDo+X+F+uEpvjEkq7nrIL0IlPqtr5qh
TYgj0rGTzHKHEgCaVhD9VDMPXu1pV6IGfW/t/xqam+BKn7bCrbYQkRef3xzacdIidGDyRXlZkz4X
TBenKymefGnXVN8RHAX72LN1kT9nCz0SmmWZMxNsHaVKQmSyMwvfpFNB7myMDV/qJAU95nmuzRRz
mrb4cOBEtSRF6zASKZcVVqMgDuRlkd8USvj//rUpeFs6br1zG/y02UVTdfriUOP7+XkAW0gXad6u
Cc//JAcORpDUnSEEPhTPMPX8M1vkSZca/nZSccuMqMALW4RTbfCZ8A/ToeSP1uxmKi0qYdmGZGSn
las6aFD1Wr5JZEMCCaLcIeepBts88zcrOpJv8nzlPDGfNiY3TNHiIgYqpK09zlvErgsBiSNopEMU
CRRlzWIjbCaEeW//JBlOhbEG3+V8RQZO79S+xbCSwL5TTMVzfVVWGeUR2g81NlFxt19EGYbdV1P3
5vprftdLyx4f4oqTSDC2UreSTYUo94wDEf1rQMDy4ho78Ovv/BOWC5q+npTIIK4RSRI65dAI0cTz
rG/NLP56rRrwoNvpqdxgKu/+hkmFp+d8BVIs3NG1STk206BOUT3lfrsSi6dd/migypeD7kTmsWnT
4n+3X7LRtKvH/wJEJB4ZZLZ1nECYxcUaZppdhk5on2//wmkyOQlHVW4S2x7ONlWzzElVlmqmaPHg
15h2/6v3LEBq2Shf2z7+DnHcPWXt2Ienq9BuRUMtJo/gJ9znn4L9ye6tqAIUDSLwgBLkFBZVBHzF
u+gEMiKbnOEyeAUOvUlLa/tXVR/2u7X8NCbbu2Rud9tc/qQvNdegyQbTa5AxDJBPYf130XzTgtsV
V24/BsDGEjUZM4yy//BHf4lUjXilLAHdIcKl8zmtnUevo5bkwz4TBLzw9PLkrPuzgyxYEZgdjuAy
wv3u3wlRjei4LcVngJRy7Nz2gtzC/WW4raP2x/Ainu2ZECuxLgXyaiieuNqXwG/By0KbfLDaFcto
FKEa4uVhMW4fRIiMbzKASVxRJYyiRnTOqDZaLP4UkOARL1Po+5ard7NuBRBjnWEB2A+A4HtkQGGH
HglnQxyKItw3Y+BIaeMeVZZCjzpBX2tzmSvhMGHx7t0Y8O4VlslSg6aIP09Wpi5VW4Qy3XU3YL58
BCgseUoPNmvbGpcANbA/lQTv2epZTJc7IHD+E21i+PbGVoKxGigGh4+mWC7LUs66GI3WwL3lg+nu
TD+I16Z9hOt8PLhJ1Bhz7DYBRGP2ZuAPt4wxkyq3xT1umZx/PkaPIpXyQ3VIqdhPI71Bz/FGFXZD
NDljwcys8WIKf66oIzjnxjBKDE2+LNKgz3XZ9OJX2/6NjPtF01Y3Nk6SfSH8EraTmSSR7nioQUVE
/Pvv0xO+FwtJZRbQ6t4xadgSeTy81OktrNe/h1VoCptHC6ZHIJ+vvYNoTfer2Uv6lfMdB1/f4MQm
oiatIugtN2iIgsOcQhacGkrsYP+AGGVyvBNxLU/oVxedofydV6ZM1CsBO+zy8keqMXxkbLLGW0N0
W909HM4SbyIdHTmVPOvLOn8RMGZQog2W1RGQYHIySfP1SXLUoDlygDMfecUDWSAf/VgKnbGR9NGM
7C4syukA6fssd/RB3YQS9D28QF69bK5gkQGFgabebZBU6uSQrFrOL6NVqUiWnbQ+BkMHmDTKRICa
H4r/knPaVDCTt0gj28O0z2MjXvBQfpDv635K+jUR6FQSoJ48OAAqcw2QmIzr1yjQlrDb5Gl7+kuD
XHGMzsZsNz7HtPxdONdoUDwFvikQSwdCN6d2F3Zcx3AueqivvsJX3IkRa2VB/Twle3YdmYYx5IPU
g3gdfZjn09qa+NSeoQiK0Oe3onbTRYobBnXeyBIxbTR2BRnEwcwSH2NEKplsbfoor5Fg2F6RNz6d
jr5SK4JjlVj5uPx90gr6B0PQ4pws5pOcq4+k7hiz6Y2MD4DVeW7QKOm4sKfooCyO9APC3IeTx6OV
j0y6MB/1q7FjHDGuSaZSpJEUJK+IJROWPUAdMo8j9X+2SdZ3E4LLz1YtFEd+EBxlgowVsmqPmmeb
n5+XvSFk1Hwwfrge6gFVVhlRsbWe2FYyAZpvnkSZRyDiMxEnek7orJe+7KW+kCxgXSeSc5/PT2tK
lM5GWVqIGyIJImugy4etxd/Ss1V/2dXic7h5nb0yPuAtQhVnOpa+mzQQvThhEZbQdq5tryypMwKc
t+fdGX758VQdSwsPZHWKA4beyJEYbNn3BxI2k2+X0zIoZJQ7n9amU580sVJzmQE40tEquuBa+JYG
ee3xzJc/9DqLPMEsQ42jV508J2XxhZ/Px30uIK7/rOZHFtghZNrKI5Eweqxol/UFBMlVaCthZJFL
7f5liAZgTsnZ0Azb2K6/WPkZSfoj0RKmy2og4qCjIniHtWjL1lW+VW5lcCgb2M5iQqY741/+Zymz
DLWra1vyX3pPl+Maz++Mlh3hiQ5+eAgGk2mpaOjThEyai4YpnickZPksBR3LRsav+/exZY7SBfRa
D27bdYnctAEM4cC76+hkMCXxkzuOCO2jYeiAKpNQRPz/nZ4uZPM1L5uR9PbDpJSctg3aGmHqnn5Y
M1VC5NbKLg15XE4OV5BPceU9nue7Mx2VX+N4dae7EpGvO1i1au+dkAzaetCmfKD4C3yUi6SMohik
uVGokUlw8boUy0RVlZqlZ6QVFf/vetzhki5KFN06QoQVSdoLfM7zuOcjyF6O5oxOZoNWfpon3+xe
00d98P3u2B1r95O0zpq+uSgKv88WqqOQGwUDiigxlzrMCzXqNaJwXWe7XF9x5B/7415JDZQjkVmh
fAaP08/T1Z+biY6IET3993u5lBVt+ayMSVbfaC6LuU+fExX4QJP7TXCUno++bc+THKcp+AKJRHao
kTXy2bg0T3ckaEB68UaL0wK3Pehz6inpj+igt9Vr6W/CQT8aWnN2gtewYkfe6WVHTH2Fr+1/d2zs
RwyJCSyW2a1D/lX61Xb3QAQiZcKFdYzTmuj9kNtZjQwrRFvh6V4EWHKWkomkD6o1MNR/XJdPJG/y
S1CFOu9/2Cidm8/w7n3pwaV/sAGvlrH5ax50UwxXkDM2UFTqU3W6FafkUlBUdlLSKVTrJGI6pBi/
10pJVdk3UhH897VIVYK8L0XKY/ch8kVzUgON41NLFXBoZITc+tzqk8cQsmQI9+svzRims3jc+d/v
jbRNYwlpU5nnIzPv6BAdGWkBvfWh50XjjiRgVAWo0K4d+eodqyUmXQbVh/TgUoZhPy3t+a0VVERl
SA2brsxSYBxaYM5vtxWbbAXAd0N48xHBzuHYZrKmXepau7eqcwyDlxsBY9QAOznzez0PxA1/aU9M
9BqWXU0fNpOBCPYijab1hP8rCxNAvqofvvEwJBkwm6qVcWzt9hzppRPKQI6tcrZQfMTIveKVEqCR
UMgIHIQF8uec50Wca4WuFmx2fMBkau1vJnUursx+1eCD1lDDLA49wzLiuu7pT3Ee7RTZkwpRNt8f
z2sJDbUuc+8efQfgyrLvLNh9c77eEF6kQemzBqRhVelCpOGh9RQpVqssmdSC9GGhO7lJpuqQf3Qe
aCbzorou4bPx/vFIWMYtUZVAWe8yrpY75LrKrAu3rehju3mJGz12zJFtAqjJgQ8/h6DYohdTVv/p
6aFz1V0b2ZLDmDglVXnUXSBUXhCpkxYp/2rzqdlStYWuGybc/zKu3zlF06/I2x31/COfxvth4sFf
NTO0llicSRcZFhO0BaEOZexISF0BQiexpyIFIDoi3V5BY2ZWxyatEeMBAC2uaW2ITdFskgrveEMk
I0XDVeTHi8XPkXYI2vIWHV0ubqXOLnZrclRKokXRaq7Alm69EuLxbkQVNlbpET1a7t8+y89Vvc7/
85hhhhSUQQE+W5r+MOjAuOCt6igIez0H1hL03aCRpI3tu/foekKa+Qrd0J8U7GTq+2prsEq6YnR6
EXOHYFOlR36N+RjDHQypk+HilHAAoW1KX0ZZpp2Ml7K/K+jj/d1/hVRhtu+RQyoqkz98Zt+LZG9W
P60NaCT91arGiARvlmit8sFydirEQldhM1L1sDsx0xz13wA+/kohX8wezYu3M+t+R5bUGzHyx/2r
Tx4B/pBvGFF0icnlQKFxeO881pL3fsht54NtfCovvT+d16xPXMdmvscINf33zZdX4eMmfiRibl8q
QDzHIzfgxZpr5eoWJZEdew9f8nH8pB0cmVP1jV0gbqMXJh+Y/yP5Lgm4iWYc5iUkrMgQXAPNRt24
lEV30TCMu5sQrGbFXBFoKQsGKgg1hNILOEpw/AxdfhRf7CnqzakFKqQb413hy7+7GATLOFtwHXE8
y3KJP8onZjcAjyWtKDhQAd9us1HzUR5XJGpFhelIFoarb0uVHcmXJZ8Rt2iRohvzCOw6a5lGdAOP
d168huZge/9yTRe+wm0u/PwftLAOetWJKeAWBEEux4imWRli0EkHYK+8CQYp0zyRHoe3pD5NsQns
54c/xnhc0I62Vm+capRmi/iGYyhQxg+EZ3GW+NJPL+GykVFNBc0RzgwTUl4Z1nqDo+dMOBazwrN6
+rPiq7R1b1U1/jnsXKSWgMh8/brYsS0kJgAfGpic/PSSDg2cdrgtqfiTAWvtaqP8sZvcmQFFpDq7
2ei5212j3i/J69zi9wpLQztfEFsyRuE3cRHN88tAubzsgOo1R1gv0Rq4fDGPp/kYhcKJ17K1u/J4
yD3kS0V2TK7AvRqmYZ//oyWRgf1RretilXpToYhlnx5DcbJ+DqX5V1w3cOHqXVFgTSlCpc2hpOaV
4YE7y55nggw5/E+ni1lY2Jm9F6AZ5Qfxp82X3OsgcqgV9g18x2Yoo0Sn0d7+9lDxcZTfxdjjy8fx
8omyrq5XKvmhYDCXuUcggvHRKzrMqTUboCscR9MN0ZOWLQ/webCwfpiKbPIvYH55bTd8ji6xslLg
5rziJL/f2eLy4Xhj2IxADyaYzlSOxFkYCDiBQ5jR4Z6BFKSXT4Hb/8nMVACOxhpF4wmXfD9o6nVa
iBv4BNwZsGd0fxgJBZU0y/WSjy78a2Wf6hpdrAhmeKa3RzAsm0VLcfgVwF8ifsKHHOfV0YkM7R83
tYwf/T5nspgu264QRJK8X1JCj5mGDxM=
`pragma protect end_protected
