`timescale 1ns / 1ps

`include "softMC.inc"

module instr_decoder #(parameter ROW_WIDTH = 15, BANK_WIDTH = 3, CS_WIDTH = 1)(
	input en,
	input[31:0] instr,
	
	output reg[ROW_WIDTH*8-1:0] dfi_address,
	output reg[BANK_WIDTH*8 - 1:0] dfi_bank,
	output reg dfi_cas_n,
	output reg[7:0] dfi_cs_n,
	output reg dfi_ras_n,
	output reg dfi_we_n,
	
	// jun ACT_n
	output reg [7:0] mc_ACT_n,
	output reg mcRdCAS,
	output reg mcWrCAS
	
);
	localparam LOW = 1'b0;
	localparam HIGH = 1'b1;
    // 6'b1 concat : jun
    localparam tmp_slot = {ROW_WIDTH*8{1'b1}};
    
    // for address loop
    integer idx;
    
    reg [2:0] addr_add;
	always@* begin
		dfi_address = {ROW_WIDTH*8{1'bx}};
		dfi_bank = {BANK_WIDTH*8{1'bx}};
		
		dfi_cas_n = HIGH;
		dfi_cs_n = {8{HIGH}};
		dfi_ras_n = HIGH;
		dfi_we_n = HIGH;
		// jun
		mc_ACT_n = {8{HIGH}};
		if(en) begin // host ���� ���� instr ���
	        addr_add = {instr[`RAS_OFFSET], instr[`CAS_OFFSET], instr[`WE_OFFSET]};
	        //dfi_address = instr[ROW_WIDTH - 1:0]; ���� addr �ڵ�
			// RAS, CAS, WE�� �߰����ִ� ���� �ƴ϶� , 0���� ä���� ������������� ������
			// SOFTMC���� ROW ADDR�� ä���� �����ִ� ���� �ƴϹǷ�
			
			dfi_we_n = instr[`WE_OFFSET];
			dfi_cas_n = instr[`CAS_OFFSET];
			dfi_ras_n = instr[`RAS_OFFSET];
			dfi_address = {{ROW_WIDTH*6{1'b1}}, {2{instr[ROW_WIDTH - 1:0]}}}; // MSB *6 ROWWIDTH��ŭ  1���� ä���, , INSTR 2�� COPY
			
			// ACT_n�� LOW�̸� row address�� ���̹Ƿ� 0���� ����.
			//dfi_address[135:128] <= ((~dfi_ras_n)&(dfi_cas_n)&(dfi_we_n)) ? {{6{1'b1}}, 2'b00}  : {6'b111111, instr[`RAS_OFFSET], instr[`RAS_OFFSET]};
			dfi_address[135:128] <= ((~dfi_ras_n)&(dfi_cas_n)&(dfi_we_n)) ? {8{1'b0}}  : {6'b111111, instr[`RAS_OFFSET], instr[`RAS_OFFSET]};
			dfi_address[127:120] <= ((~dfi_ras_n)&(dfi_cas_n)&(dfi_we_n)) ? {8{1'b0}}  : {6'b111111, instr[`CAS_OFFSET], instr[`CAS_OFFSET]};
			dfi_address[119:112] <= ((~dfi_ras_n)&(dfi_cas_n)&(dfi_we_n)) ? {8{1'b0}}  : {6'b111111, instr[`WE_OFFSET], instr[`WE_OFFSET]};
			
			//dfi_address[111:0] <= 1;
			//dfi_address[(idx+1)* 8] = {6'b000000, instr[idx], instr[idx]};
			for(idx = 0; idx < ROW_WIDTH - 3; idx = idx + 1)begin
			  //dfi_address[(idx+1)*8 +:6] = 6'b000000;
  
			  dfi_address[(idx+1)* 8-1] = 1'b0;
			  dfi_address[(idx+1)* 8-2] = 1'b0;
			  dfi_address[(idx+1)* 8-3] = 1'b0;
			  dfi_address[(idx+1)* 8-4] = 1'b0;
			  dfi_address[(idx+1)* 8-5] = 1'b0;
			  dfi_address[(idx+1)* 8-6] = 1'b0;
			  dfi_address[(idx+1)* 8-7] = instr[idx];
			  dfi_address[(idx+1)* 8-8] = instr[idx];
			end
			
			dfi_bank = {{BANK_WIDTH*6{1'b1}}, instr[`ROW_OFFSET +: BANK_WIDTH],instr[`ROW_OFFSET +: BANK_WIDTH]}; // MSB *6 BANKWIDTH��ŭ 1���� ä���, INSTR 2�� COPY
			
			
			// bg, TOP���� LST 2bit 0���� TIE �صξ��� 
			// odt "instr_dispatcher"���� assign	
			// jun L H H -> ACT_n => LOW
			// act
			mc_ACT_n = ((~dfi_ras_n)&(dfi_cas_n)&(dfi_we_n)) ? 8'b11111100 : 8'b11111111;
			
			//jun : RdCAS, WrCAS
			mcRdCAS = ((dfi_ras_n)&(~dfi_cas_n)&(dfi_we_n)) ? 1'b1 : 1'b0;
			mcWrCAS = ((dfi_ras_n)&(~dfi_cas_n)&(~dfi_we_n)) ? 1'b1 : 1'b0;
			
			dfi_cs_n = {{6{1'b1}},instr[`CS_OFFSET +: CS_WIDTH] ,instr[`CS_OFFSET +: CS_WIDTH]}; // MSB 6BIT 1�� ä���, INSTR 2�� COPY
		end //en
	end
endmodule
