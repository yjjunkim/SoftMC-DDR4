`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "XILINX"
`pragma protect encrypt_agent_info = "Xilinx Encryption Tool 2020.2"
`pragma protect key_keyowner = "Cadence Design Systems.", key_keyname = "cds_rsa_key", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`pragma protect key_block
C0oJF2SuMa6l5UTKL3oQ8NzIzSt0InrgoMNkISrJfbH+L4MIoyjcJGHLfWlSoL8sgNnJJnewfJpv
YfYxDbNsYw==

`pragma protect key_keyowner = "Synopsys", key_keyname = "SNPS-VCS-RSA-2", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`pragma protect key_block
T73gREUbEeEcadgcm0Fok6jWAkVLLIAj0g8M1ElpcxW4VzJb7Eg2z1clk1vvjr+ennzWkPDdCqSR
7g1wInRiACjYhCUiSW+M3ZYhyRrZqbojKW6+M6XtNNyn9fcoc4CNqjb1z0dKzQN2Ed5VjTvH1b3k
XUlVT3178PUueN/MvG8=

`pragma protect key_keyowner = "Aldec", key_keyname = "ALDEC15_001", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`pragma protect key_block
Zp3QCPiy/URa5u3qn57TB9bhSAk9uQ0biVaxe4uWXuJ7pemvtklJ69FjvHdb5FlPJdQntbtpj0/f
edX5k/wcAwuTS7H7DPI0Ws1Bqz6CKOD4xaTHv2oslshZRaRQvIrmdN4Rw/5qp2ZSG06Xi1hSxVvK
Jg0eu8PcJGqYXLYgb5QC7INxxreeqds+4xrIlpd1HK3jxui3Whj9er/dQnJZ+TMX0wEAQBixOsBG
gnogY/28/lCm/qKY5uKuvCtCyYlW7kpiaqwLtVfSOPUBakWeQunH87r+ZPutRUEJSHSqQNJG7+4t
N3FqL8iQR3HwsFNLhMXnNGbvWTOug7VJ8JNqTQ==

`pragma protect key_keyowner = "ATRENTA", key_keyname = "ATR-SG-2015-RSA-3", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`pragma protect key_block
WlpHIH6+59sUqAlQSWev+VnSCbtuwXM7bkHr4rCUbCJtTzC2OvCApSZHHGXFjCeg/5bXtIcJ+Z6g
fgSBcRGjcyg06GJjida88LkRfX1zal7u1LQZ/b6AKUY6GJXA8fgPa16oGYoXZCRglkTA0usTHpvU
7zVrw1GSAcV1Rqk2JMMs/7odJmb3bPnHsmAPM7GmZmff/DMbNQTrS2NWKvl6Y68UbMLeI/+wL6n/
tED2pvdOQm6tYXELI+YSUhIVfyK/Rcy3S1S8Nqa8E/034z15I/GKyVdJpVb6rX0V+sIfvzBHjNBp
v5XcsEe+J5UR6CR5b+OuhKT8AVnqMVmm2lrdHQ==

`pragma protect key_keyowner = "Mentor Graphics Corporation", key_keyname = "MGC-VELOCE-RSA", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`pragma protect key_block
s1auGT8s07pA5X1CC1iqJE3xKUF37HebCmECcARl84x+0IqQT4kdboNEDw+7/H6a6MdaMRGhTeef
X922orJDDURsbC8Xt2TrwldYajGk8jNMzNqfIuVWMLvijNTGfyPl4kUyXOri6Y/HpCMAiqQTUn/0
C7m1aWIFJDiPm2SuNr8=

`pragma protect key_keyowner = "Mentor Graphics Corporation", key_keyname = "MGC-VERIF-SIM-RSA-2", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`pragma protect key_block
Ei7FxD+k4QZBqit678M6N0vzExc2reWl5rdBjfOMq2fMZ/ljOAmwMn+uaUXPYEQMXm+/5admVo2G
/C2zPOsusl+osaeETBe+bh8KF27lPvYzGK4ziQR3Hi3I30oOyo4V9GjRSEZz7reDE2SNeUnB8RVz
B3g93eF5IwwjnW2AwNtgf6E4gvYQeRoPk9UAN0duY/fH60P0Wx3FUEcN5sey/ExJ3MmU7VCZH9/v
U/6Wj0BdwAleZFNFfBxNyQHnVS/wE35qsyb1cOonZu/fsEMcbav/p03XIvoRmdl0X5cZt8RcQdav
ojYJeAb/sCrZOqzm0FpR5M4Owh4aRCCj/kNbrw==

`pragma protect key_keyowner = "Real Intent", key_keyname = "RI-RSA-KEY-1", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`pragma protect key_block
wY9QtmtV84Now9Kq9cA7AwRQ7O4mNcEX8FDE3uCBJzno/JF7N3J321QnQ0dxXW/iXhyYnlCuC2Va
oOnDA5SidFCVZ9Q7gmc5vUg0fph8Wng5BwwPJ8XUP1mHqYKHs8vYtA9G4lSTuUBj9jRhLQQkf3TV
IE1yzmILHl/aUpBqmkjJ6mRZo8dQS2i4Yc9NH6BTPRQDS0yFgh8/mexim1nT6vgTgNf14h7omDPI
amNp3Aafutw6k/xU8eqYRWR7pytlYHCia7+HHjwBI7dUl7T4UjmG1q3x87TmcZ1q2u9vHJsEIMMV
34EVPExsKjtifd6Dd5mguDr8rIKSaRCF2tjtkw==

`pragma protect key_keyowner = "Metrics Technologies Inc.", key_keyname = "DSim", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`pragma protect key_block
eVM+E5yFaaEW0df0uVjFsuziATF5vfG4cSmmBEuGSLcO7WzDsopPqRvwLQ/P2P+nqdPLXPj7At7t
U0/Uoeb8h2mikT0Y3O4xYwsot79/uJ/fh4wLf0kCYLBvH8+4eGdt+OZbMATC8w3MMDU/Ztey+dWx
VXf8/lyxU6R/Y2RF1AU6lGpB/rar5mImrHV90febD3ItbvH1TmTnj8NJDMO8jvm4xuUtJojg0Nmj
43DvyUbmQCOK+8gCjCOyQhPMdTh5p+mx8x6fIuHL935kMkcogRtUZp/3Xp6dlMP35OJpsEogX209
xaOi6daJVsalpJOhvKwOEwRsC1uQD7w/BNt/KQ==

`pragma protect key_keyowner = "Xilinx", key_keyname = "xilinxt_2020_08", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`pragma protect key_block
RPpz5aiA1FU3P+Y4nj5b2duqFntW7YLQveNMMRIIbWzptbnClOymdlEWJll+G1/aDsYWhqtwulkx
/ZfVvXbuYhuDIgOmOQTYxBkrYPxDN9SIGBuyZAN8s9OShmCUJ5cNv+nog+9fJ6Bvh3UTbZ2IPT7Q
I4tpfDJnw8MlFrTEULEYa4JuAe4NHW9lwZI9FVlNY/53wP8EYxF8OJmPPts7wQSzH7XnVytpXV+p
wZ4L0VtXEvZSCC+7AAftazTSHzxX2p6FbWl55UOIHXC+rxevOa+eATCnR8PO0GwNB5VyH6IhvH04
f4ifslvamlFYShLgBLBEOjfwmCe/0MdAwDeQ7A==

`pragma protect data_method = "AES128-CBC"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 15104)
`pragma protect data_block
SqC3s74hTjR+1MFnTJCcueRiGlzqJFhYh6eWPKALuL7KYy2lbYdsr/9zqMa/25XHfuvUp4fSvxcF
eSSe5S8ZPx7owrOIEftAknToJrUrCvFHgTL2Sxzf+Fqaig6njBgc5WncdUBRLvinZ73TxncwfXdV
37ptzKiPmOnRJtbCnJZBcv5HVBtpFt3z9hn1d4o7C68QEAnYcRX3LjyqADmWwIfQN9ek7/3CPPVO
g4BMvmkJ+11pqyuBHboVaat1/VoaSGWIOMxCIKeFmKxNo2zTWcURm+mRIE9yaWSQx0MKYKOdQL0Z
FN2/v4WI7zD+YMPorOaoPt7ABhgaj6bZrQGVi8bf6wuUo/JTCzZg3r/rOyMsLjN1rGXTh0Nv4Gtu
kUrk6tbTqnR4LkM+9MTu5MYRlhrrXgcXFffPpAx0Q3b/2c0tOwXmvZCkaF/Gz4CIdAG4A9wbwvbk
mDp7AHKcLMOk9Nc+iFdITwaeS3p5SwlwT+9e12zsOTMee1jieNG4pV7kixAkA8p8bBLTP6y5p6S0
pfCYHDwghu7Eje2a351anog5Uy8OOLD4ioXQOn8NjXI44U1Z7+lhfHPdWJMxAiu/k/r++eBGxzFh
4138qODNq8tO3ZuAy4hK/4eEfyFcvEZwjF3Hb0qyhvaamWLYBHcE8sgdRRDgRjTH6fr4LGudRoC8
cNYsvhRKyrTy0nsGQIzlYcG8eA8oMtr76ZAGnvvgNfMK+DOTNTppRJa36cGpJt0aCIZEGEYtq3qL
ly+UrIe2kkp6ouDASCUlrgva5dfzkOcB4MFYYtxwnRt7fJCfOS9wWYpl1JoibTxB7JhHulutFQ/L
YYIgaEuDU6ac0DBgK/z7PIWOKmVAs1Dc3Xb0J7qDJn4srcEgeVqawxjaZ1HBp+xN0F+3p65X/JJb
o7/I86EiCdYD6ONRKFzOXYF5vMVXkh+wc9mInUCOk8Ueqvoi229AYXaZHsK0EJ4mwrb+0aKFWT/Q
shYNhq27zAqiJkDhtdsWrW1PAsE+i7w8ZrRYmGYspDn2h9onfmnDN3urLYyHGOQeiyoQ8hYSeF0O
WfdQlCo/Ds5zOE9qoGysUM6kxeoIs9HrbbJVv4HtlVjufjbp3wOWUcLJlKnaluSIzloCrfgPaXj/
aCHOMZUEwI+BBoVWRXJLR858adX7RNLTBZBdB31FT+HNKLj+3V5+T9ArKvM+PiTKuHNO/Er0U+4X
hEkdMPmZ5nZkZE/ttmR7GJbAaVEVamvz3kZia8ZplNg4EWsXuzZL3QYd2SA6gh8lQp91o7bCvwHX
dk3g2FKfyJW9QGnEWlnRTU+vs6gahYfYp6Ozat/lADW91RuSWmA1HoC9iZJv9lun6sOvGSZEjxaa
zOgPBoM5lRZjYhxjXXV3j5VHoCXt5BpzPUHw2+GIKwKOPqWwrGVzKbGGyZYo4T4RXvsFzg0ZsOHp
ZwPscc7QMeYSBU6dsaa2kxCH0rNATSjf6qIlML7xBIGo8X5ErAOyo1hH/ZQB7clCJZnaxFqDHCVp
IJFBB4VCksazkv89JvQzwvbtjVjmc/qk5At5EfWKLzVE62oi0W8z3yFdM25aU3gCkMTDKVn07xS5
m2d0DdFdEdhk3ylRgRqQd0+em788o23O+NLG8/mxUQ+XAXmFIrnam2zXZlAHr59xY0cWVfz+b7AS
P1vxrnDeRwUTqzUk7+TOHddtvYmSLU+fDK7treOItgmzsYhmJgHpgv224Ew2ImoUxuqG7Ad//OcO
DPGH/oii20NyEwV9xfva9fdudvBsmZ3nGEuSOWVDTJt9QYE4TdliAofVmSnqii2gYTNV0CHVFLF2
TGkF6BxR+VBxpISk5Da6+5TJaQV1qnswwfqzlCk6i37+VXKQKs9k8HGtoyXSNbh2SskLxe7Lp/Qi
OSHvdkzPp9n5cCKabXlz6S9HpQIlQhM0bszn9tng5qTD0XyfsOFdT8NWjVQ8ytORIq9Kj1b1lIeJ
wXkXcj8DKC9OY5sMMko2mk/Ino/h/M4htOMm+LNlZfU62zS3Jq6JXBJxtwEFun1xdTTA6NXCKrqt
j9kBSS30ba9gLQYFQ44S/6/J0YRNnFNitz4pGq13MrxSIWxeeUHzZ8SFWuo65XP4hs4vPrMpw5j2
SOzEx+syMHmxo7FslpJjijJDlXH9pP47BpL7p+Kr6ahejZTA3Fd/BJ9MWDFv6ocV4OA4fzvZUo5O
+FpbqOpwWw1hNwCVWiNbF0uv2u56nDtbeyE2g7QkEAxim3ZemZ7teTpoMSekNOTz1E6Kx6R2aNCQ
3UeX1n6KymbEfTf8pa2j+F0OD4S7aAJX5sXWMytE1XL6zISFjqNd4c49E8AV9IMcKNQtPtNJ0sVv
8UYjmDtz53EvJr3V9/F5twUPshi6YOCLEN2w8b88rVgzi5VnN5OGOXBg/YZbZB3QBwzgYeFX3Q5s
k+kjQoc2qhXiazo8W3JaE+Ch3GmFgH+UqYWrKAeVWwtUMXU8k2+/G9fQBSWN8TUfuAGyYXdPW6o2
gxBKif0tvsOJGddSivV4zAxUC9wNBaXI9/460GjYqAx2AOdL4F/xz2o1CQ90oUSfFIG2yet7+QXw
PS30cvqr3JsfpZFXvaJfF9CWlOiT7h7/uQ9lQkGmLSC5R0cJ9MLmWZ30hIYAKMmLe30bcMnJ3fWs
eNRwO2kTznGIdhw3sr62qWU/h6oHqsxfnZdcHtD3iDcXfhu4SAYzPwR8WsnXJzj5BFAeVTWoYYOm
rPijQu4PxNmXh/krbs0lbAXaxXJDN55yAqE03RiWrPafpiaU3ww2mRKE2NvRfNPfQPm/98EnvN2w
073UCjVsDNhe3H4R6dEZBuMPi+KZnpc5TOOuy5PYCEHkZd91W7Rp2IVG8MwQJ24aEXYthca4vAQ0
HrmSh12Eb7GDk7QxFtCZLJY8sKSHcuQB8LcbIjzFjxqYItsAXnUsRguNpxeBOTPUfT8wk7hGJUuA
8R+/qFycADxlddAsgWv4/K08fSI1i0SYGdOJb9SjW79k3YqT0j5pkMsjclorjI/XmnyRAu/q1k/o
XqK/+GC/9B+thTimz7BKobHgRzeBKUumvrUyFgfD1lzzob/O1YejYGOHS+eYkhxZrG6NHCNFO7ua
cSgtczWTgUZwgL9w2WAH7R3SJL+bnnGi7rtUpMcWsdzeIEuonGiJ0uj4rkW70/2CLu8XUavL7ykR
VsAL9eQU2JFaxztstFufFU5MsBVeDdJx9TLEo4Vzsl863XQYrZJFa9numhZYhUsGJYpRYqtHG+kB
WDEeBjnwmoFmbY6vm1TXJvNYimiX73Bl/g5BO+p+yzPEIdTl5z5gDO45w1XlsQSlQvzSFxxwu77l
23mItrbvyKWJU4o5Y0FKBJdWBSA13D/WiSXrZ8nUMQevOQS4oa9x467I7s9yfM/hFuOfsE8VsVft
8FmOXzjQ/jQb2YcC5gWml3IMzeE72xE4YNZpSAVDCD6BlrwUlfmr/z8F3pUc46QlI3sVekxo7EvE
zmv1ezDnDznFV1da2FgQ3873UFhAdj562hyISjTvaMq8an9uX4M9QwFVqJaSDDFMa8SBnnTTwk7G
V3OA8Jc4Dsf4BdUt5oLuCoMnC138ijrph3Q8lausGEAqgYx6ghxmMgVEy4ImcY6AUUXuqnjOS3sW
6GoDUB1Lxsbk1+2A9mJHRqKGPsuK2PFMihOMYG90ECkM2ufOD4/6NSuEVt8ZvRa8D7LfHooHcEf1
9at8Y3xY1VbHuGBpoRqXc/rqKQN4VPywaZDF/lOOGhC6PpMHLuhZGk99IfYmUee5g85oUT3GnEhK
AVuxBcgkLKAX8jtwpHVfL6r2e4io4DXmihMNq7u7BY6OaZNuXqGUvlkhDam83P7Yg6KInIkBigmU
yf+LXNXwcbd+6jJrgwPZqIvugOAPXwk1zpduHDd+tfllNZ2wpRS1ugsY63PceBtzvp5P0f9ejomj
n2Ks+5ZPhIra9ZQ5J9qGDhVo5IcP6fZG+/Xai6XWb9TxjZJ5i9TxTZyHMiWdxYwnZ14svkiVB+8V
Tue9VxM8tJ9jREphmqCtPopzwTyI5HISwYkUJz/WdnjKBRjykAKpU933vKwE/EDFKt2b335FZhXn
D99TBgYy5nj6G3yKD6FQ3oxp/P+iBI5VZmf+NZZ4KldQzG9d7h9sWVQ9TSz/9gMFes86cnrJdZx+
0zchXyofV8wdpXkzmTnQTm3Tb3tnXGXnBcsN0/K5fPDNIr6czb4q8kZVhf14Xd5fjcyB+hqCYLnQ
nrhX0OJAj2mjrb/iD5BjOHxjDmzC/Qf61aNWlUdSXXKy7DhzYgJi274SUprI77AtXxbP1G7ZKrxU
VdBvSGyYMeebZ65cx5r77NhkHL+BH9OsUK3UYJUhLyr455ktslEM+gHx54LefGOVZI4W8ecOSkyx
mlRUhQ37DFRfxZMtyFbP91K+tlv619+zNi1+F7T5+/F5ypcvGD6c8uKC7XzvOzVGXYh7lSyNvUxX
39qYE0RDUQe+a/b26Sh3x+NMAqHVKIawISSsNWsdGN81dDDWw9OOKLeWryWn16K5BLkTL7yB6SV3
N1yV33hU9H3qf/Lgq/AD5NOEVbipnuqJAW24Btq8g3qKj0zi3RnU0z5FjIu6I60oGaBRCm+oerxx
QN634FkGyDicL8HfZRbCAck7vnyHdIljlTtTbZ4Lw/ccc6eZUXKmrilRTjhkxAct5Z2hSRiwersp
TBn/IZf3nSdVePFadCLjuYOjV97q58+qWLjL9LQlhESGcMETnyChqfF8zj1IAx3w9rd3xFYorr89
pB0ouWXU7C6O3S2xsUR6NAJXdX0WEKKOrCgHekuYN0BrPyMtF/IUEssKMLjCf7hfizrKdAC6R49D
P9fTgYqZZv0M3cJ8m5e2s+u2i7r4tjlZWFEKkqGtDQVaGvoGfk4uNPCmtKboqIGKdZULoXwxKPXJ
zjWzWWwNVbuCrwRqrxLBC9ImJ8n+Td94YMFIrdTOGAedY6xzDtfDEdpLHTF+C0V8C/ykvDlhnJHg
xfG02xFsaIyvNU0sjMXKlDEcarkl1vYIZn2aYvy4Zx3W5AI6fmXW+EfqWltkvp19P778iByf3jXp
p2Ns/SLue0P5QND6SgT25oDC7uEUQspy6um5TbkDQ6Wt26hryrqtyRl+TUmQs61vhI6sqeOtWJiP
iTGVp9RcQDXiAyllE4V6DSmToFiwQVqwX0v33ZaoAxLRK8wEruT3u/X3hrb+b3ZJJuPLmW5SEPko
LQZEMGsAGbmK7TWbqDzPXsYY1+Y6VI9SX0Cm0sRPgCQnsdFOz7+hMW8rg9cfK/XKuZFngP7T7x6Q
YUWFcK9NWa+/erxDQ4c5aDzxPNjBjPcdFMt+7oavjvqr52gHJE/69XZPZZxeVZ+1thSNT4V/Z3cl
/iCxVlrVDAEdE6jUEZzYk6GqlEXnHTCCIaH3ssMKtg/uhpwvU0SbFfEAd6cHg4YP86vG+XrDKkeR
o0/LdFXdfinWFc2pMc96ViXCohPlYQEg15eSoKVe3NbGI+FMQux7MoAzDeZeD96YYT3ngWKOsOjh
H7eHtco4l9MuEetsusm/jgx3CoDOPzHaS2oiPTYIicNbFjjITReNf/CD5O1KlZkv2BQQNhzqMujv
UGcmqSTzIbinCWTWKVKC9wJPuG0dpXuhLlTKI/XtzaylPqHj7mswCTe2Q/U+arMgr78wJy4Lkvk1
9YI+05n48+/qD5oJzJ2nvxbO3OUDz14B1AM+X0u6EaYp2hAcFY2SeHs2CPlhdCzItyZfVt9hrqAF
yRHJdTvEzl39la2OvJRcoEjetE+b5Fny9bo8NjCQH+BxHyQx4OLAFVrkQzPgR4tpVL4OcYD9uhxF
b5DdN/sAl3wkBwCKLMv6YmaoAqPitzQUEyS3BiRSNAVnl1a/yVfFfmAyrhJgk+b4wZTfu50z/+As
Ac5eq5am7XljSpGCvfXlYemz3JDJ2ob3+OUymsw08Yd0zi5Uvx1jbtNbY71YtWyVQmcw6QRSOcmV
2/kw7GFvWZtVkv9I6oFGN/PbeH1ikPeuD9OgeQaDwMLZdEjtZC8YrMKXc3rPbRjC/Rg7+yw6+qKW
nWgIeLFVdLEnfvl0HjRhDEHi6IAAJwg3lxVaAS+wN/mB2vcLnmmCsdpgyPslEKIZbSfk48kZpXwI
SMUhZXOJKJQ8pUnAIQ35eVkrD9fN/H3Gon3y3a5LZDsf+SBSMkcdaA5AsDqlI3rDtKM45G27CWIO
tpSwQx6a57syuIzp2/8lnWOk/LSaQdN26TOm2NG1zidONi1PRMfLlMc/tXSiPoCWfnw5p5sAixBe
n7zvOpFiUEUp0GO5YkxDFN4MBg5q4x1isOADToNYGBy+4UODVZafNzigDKIdJx0tOAs9NR/EZ1Wa
GglS9Ku/dUr94GCOqLaB8zA09dSXiaWhVUb/e7nx1s7eAIZCeE368m9YyAINCdHOw57V0X7mFdQ0
/u+ymn7Ss7CmWHdbZrH4aUf7x4TBqrlUhKQMCg6AOn6bsyFFzzz9BdyTBJ0dhkGUWJhhOhnQ6EIf
/sVUlKEiKC7DTiFqJG6I2Dqn5HRQSQ/UHd5/ilazBkjw+wFjOm+gmbwYTUpxx/UGwtXZRNgsl29Z
0edKCxH3bcLwwvdliq4VdHGngAAOzQ52XlIZXMAuobbGJQPJNDxy1KFIe2Jw2Q57RxZtpCCdP1/r
CBSZ0drr6Mv7N0TdO8YKqvWHV9ZMFYYUmPgsY2uXoiaxkcrPjRX02OtRsFHORI2/MYghozLPEsL4
HdHXlcjlcLq6SJUQ+j2mTu8c5SrbM+rjuRVQo1GdGKlwweqZZOBNt6Cr0tQLm05s2qf/kUs6pH3+
+Hj4EboPBjui+fxAleqBUqmjaVE7OJM7At8uhHAOv4YUxPexktyEG5Q+IwK32aaY0wdgP8xXS6jx
HRMI075YXz4f9vW7DHRcTUrer9vyx6i07bw/1dGTL8DZYBAsF8ESBJWTQGAY4q+pAfY5kDm7ssza
nncF/wgmP9L0Hn/vz6G6iLEfqLJnXgjPMN+Ty6HA5xFYVzuJBnvAciKd/vMZbuQeuuGB7XqCotc8
EtY2aEM5kdFTduuf3bFaDWaaZioE0O/MmeSucCe/2LwmZrmCwhOxYKWXZRdN/SbK2GH0IzrtT2DS
daf3k4tfjoJ+U2wLxoaJGN3DsUz4SMqezIGCkGe/QHmpKoIxa7d7UFo59YLzEZ5CedBx5yB1qFIF
GHFJf9tF13bMhchaT/FMcclFy0R7jYH64jBVPQy/hN4eSus1HC8673oTmFOud5sQjfKNXQ1NudrN
y+YQrCZguqXtOQtEyNCUuMnL8KwgGKUzw1dIfdaL0olAjqS6cpeGcNG0d2+SQV0jLn3ZQWJcPEW7
DOhoIHSb/ggT2oMJfvrPXQ+VByJTctP4laG0X6l1t5HuQmxwXDCO04ug7eK17nlEc6fxmVlGffKa
tZBB7+YnNW/kIiIXuBCp3w/4bsn1P7XcKq25zxZkzrLZX/XOfXJBauY1WIcb3Maz9q60vaeEaSjQ
/2OqY+Nk/+5/LASbS8D9MuQ7HONWFw9E4FZm0aICJb0zE31hdNCW6vB+qdzr/LpMIhQVJnfg77I4
nZJkBiocSso9ZH2l0R0bLBPHs8K3OLm0Mgz0+yfeZXVtxb0TAdVt/ok44z2ICZWyJHEbhLBvXArV
ZFMuri4KoxbEBKMRWSm32tZDEb7s45uc9db3r/pa2jELxatm1Q1h6lcdchB79oLDaKUohuNEY/zL
iZ9PGFva8BeaD/oDltU7x6BWqZZ7vPaR8uRZCy2GqVYBZm/DszakDaDlDc7QvGyfBl8HScAz1Rjz
q7nmzz0jpVam9QUSwTAJgjco5BlgAQ4HyIiVajQfzVvMUsl13ocomPs+bvHOjn3QDf7BTVV8fqcV
wpI52SmreLHEl9vBiCMPo38VSmiol3+p/KeLt0diOMCk6HYLil/4AwI5E6fgFmOymHfAxjrxKZ/s
OX22bnH9QHuD1SGSzbKmsrDc+u3B02K7uSkFjX4Pm696LwHIni4WuMBXS7gHwXExHWMaovCq0RjK
BeJURJWX+BnDkAcRhtFnoUMR/oA0yOTPa0aW+dUzj+yCqAl91ccGLiYOlk2inTnLb1K0RInoMcKn
ReNP6d+AC8P2nPTKKVh5lVb7oYnnobs/Xm5j6GLbDwP1rP3kWt+6iB2kRq90OtVuuMKyk+Hct3/b
oIkDuTjI1HUAcPUxG0ydLZXdWdKQt1/3Iz1uLCTV5taW9jtAimyGFikrnKjY2ZsEkaSwHN6u1wRV
7ZWus2WaMBfm+WtItdh4iGJB3vj8x3Bb8/u8Kbadsw8wI3TT6qAeS5O+kLukHTPSqYks118+yY1V
bUM5FJh0Tgvu8XLEUD6xf3ltLGIctvYo1UNLKPJmK/xo7mBRePEV4jETwBy+JuhCz+RGhkXfMaJY
Vi8D7P5LsrrEllO5o1I7V6b7BKgHzZmssF+TUmF0eK+6p/gYBeudTqm3C889ybR1wff62M5qcXlQ
tl5wRgUiYyc+a6e9+zIgPig3WGX6k8Ysi15zSnggsMbWnPt4Zeb3Dj0B/0VDs9jG/XKn+Ku0asIK
br5ZYA0I8KAaVvL3HCUdD8jeDgaHb07idmN5pykg7UhLXIMI7xPBV9K8D1myL4bYn2gKR1z/dMeX
fEwl8Sv1KqmJU7MySvYqL0h4eGwiz4fj+hWnWOlfBeg10PyHfspQcaj4VvkOfNzEjJiQvQR1xpTT
GLFcVajYO+hLteo/qkAAgiYxDD66A8ujWtEJdwkFth5gTBthT+20wzGEln3h8jYE/bCMjgkwZdDb
G41MsB4MRj6tZOBDBfl79o8lRJmYsTVGPb2aKcXrvwUT95tAY4X8Dhk2fphKTaZg3KBqOZSuZrB5
OB0a52BbBEDI/IpHjEAbwbvprWd9+Qk+zvVWbN7hpXpfUbckyp4B9K+bZTisRigDL7NNxb0h2OC4
frXqtyRUp7kaCMhc7qvmdwgyJ8IHx/dPfZbCcnW7/93tqjIGCDMFlAAUzN43q2lAF1g6DCZxK58D
SSbPivsWgQzhjSpl5G4U7r/9bxiZFeU6kpD/L0owRAs4D+Jv2FW2BMY4TBc3dPYOvBofVToXTWdl
Mi6CFcVmj8GyrZntUhcUPV3YkSO80BYpRNh/fGzGPJrOTtgEkUfFqtjimFPb5aNM1DvSeDxqV//v
WciQykJ4Wh4PjRXqPR12eJ6eRjj72XKRmZgXd7dSqidmLIMvXzErohr5lVSEvWnQHo/L4tDlDX8U
uyCngM3xs4V77dDkd0raax2rMyyHuViI7uzQ4d8wPP+KCp2WoMIZOuQDTYidyXJpy8YdaqKJFyKl
8mXcKpHhfmNsd9iOtzTzXHRu0rUjco2GyyyKS2xCanXiQuaEri2Qe4MiCGh0pW6Z0xlLHQ7l+2Po
0LN0J4z8YzxVLHt0s+2F+o2pRe//M7l5XcEMUYKAKciskJuJ0ZPaLyJPVEqxKmrqbz5WEVvx762b
aTRYmRXa5w4fqATfO+ZHPyivBnieccZCjSNS+l9wD2sYyuM/vAZcIUcIrGhU3CoPKZzO+dKDQA3B
4REPNrmJ55jxEXzJRB+pjnKmW3ONX4bl8SJVNSB2WJKB9bfR+eTzvWYY1VvKE5BdgyrMUxPe7k40
J/x+2sTGPt6fxEGVyQ5RloF75FLL1VsgJgGNN+M0CGP0KkWZhQ4sFyJAajFNiB7x9S326I1CQGVQ
6d8l3uL4Ly16Le9ebL8VKKransDXletwdy0IWRFubT/OwZnE2agaCmkewkAVNeEM+14nH3BOuMvz
zT7DWNTERcY0yjaqVy+E8JXdIzCTwqclfIYkeVpLfsXAh0vUmuM66a1Yxvh9oLky8q3EFXtBuMcv
v1HGniGSEI2jTAKQJD4RZxj4FBDiu0l5W3ffmLnRMbIGNMuMAIPAN8Pq4KY9CXqsqvImBYRLiyUM
jS34kGFJH/Sm1174PY4Y60nOsABlpNXUx4lqM2/snlcxIxgJJW+kWihBg34s7UZwilEMTGYQJtar
fhPXCg7w/01IRHEyUc3qODPU0lvQc/msrvh7+siX1UucnqH7s4vHKKqrpXqG2CHhvtbq649CusUK
b5a9qObsUpF+oY41ZcsGOEsuT4LGPWj+LZMtv27KT0wUNmUCFFMyX2AilhLkGvr8wtmF3x/gfnl4
esTVATEmhnmKOqJGm6kfrq/rGlzjh/kKZlikvcBfFJDm5ohk+mPPnmA9l6Y44yShhmslLnLsrICb
jqLKU1VDWQL6oXbh1pg9UKmZyb/OBCbI7NRYZEeVFli2aYfB+S47BaZALC7y46q56/sT0dxr/0it
GftGuoHSmNZJKpsnzfW83b+qBRxFxFqRW7otHeb2QqII76KWc9rz6ZoPCT9my7YwyYylknRYOB9v
1D128w+VLQFGeY9Ws+lkzYfQSRO/t9W2jIxuVcesKxvDGeCM5wWVa9Zqjl/oWt+A8PpOYHOQUDoM
anr8Rd1PJ2yqKvKpDoZCdA9W9ONuE62KIeOOjQHsaJmO9eXXKXB6BByF12PY9CjKxwLE6f3Gyv0c
W3lF6hn4aI98cQaeDqj/MJYBbEa9DClILEDopZcy1jA67yqcH2zEBN6s0CpHJpYaFjCS4CkNrCIR
2nQnVJTKbDQ5H222S/K/vpEqcRV5j0Gu7eWN97pHcE5qnyxyauQfy9gywLaSRJsOcH8CL48FxKuF
z6VSYQ/C0A+lsbrSLAxfdy4fQSsh0h9K3zXpWlMjMvOl6hSbPtAVLgfmFc1eZ4M2f/YSF/6fm6A1
7L8jodKu2w5/6W4zQfLkpU+PQ8k+vT8DSvYCVn0XHvRDINr6SPvlg89QxAYU4DNu8TdhAqQexnlc
twhK/2DEKdEa6ONMGmq5odDXetY8clq/sRFB6ocjpyw69FtaoGI1o52EZTi9XBmm/nnIVNPeEfpo
0tf3PbZLSMk9FEzAaAUQwhLk9OHViltpi07CUQ8vGntNviw68SFixyUG6dXDbNyBV0ESOOXL6+Mh
Vm1RoeBFRSv2ECzFt6o8H3vt8NSKqR22TZkd+WkO5d8qaLsBi88N7lcFeWW0NJgpeHZWZ29ZwQkz
+q2XZ2FESe2gg3fSMW7Q32bV5ZICzPTQHJNds+yDUlH2ls/DT1CCMz/POGZgP57I4VkEiRsF/XJQ
1iHbeUEilUAVj4mb33eA1sROoHQcYrsAxoeOu5ME7H03cwNCXH+nuIjmoZ57eF14DLlJjMGFbCwp
hTzNqVn+Cqhgq7LsK0l1zgb4uurgJBvchL2QkXLsEfWKHx4ar1iLj1xvbs3WsXQpbmDEvsZb4TtD
qYxYdFQglL4/cRG4ni9UWzkn2cOLgBYsMyaW6XZcOWVMOwapw3jS4uKfOJaeUU+Yq/95eXCRUZgL
Ko2Ep7m4ZtQ1VIKqMxxJ/wgf754ZlwTdMRtsPqaaErHjVjGs/q/MhBhncCz0FN+SWAFhatOaeIfF
jjosYqYqWf522VB3KeujReBbvbCDEQDguxcvYyg8QfbGFJb2QmgSDugxFvQ60XNc51hnwicM91MA
Ue5Ggk/DQmzTIz7p5v5YWCAz4JQd6Mqmx0LcuQs0IQ2BxjNPjBRSiUmF4le9Rp6AD807ysA9Tc1o
Ggdmb/jVByVX6i5R/ryLSxt/LlSE2RRJafddvV5Z/XmMgys81Vj0LOsHvfGnULkN++1GRMwp1gSM
qHWkjReXZXDPzfTy4GmEKRr8C3LTNCkpROAXQU9gUoglpuymSE4czSbSmfd1L+rOoPOOmDXZBrub
+WSt2foHw9m3Rv+8EUboeMHrQCHYb9hvTEZtvPKkfrrVh9veyOQtPnIgIadUsz75JPAXzglXiMX7
iDZBWfLxwI68OVzVFjnDzkrcFsF7f4B9Qvl74o5i/jbXnMmrhdgJ4F9I5BodWZiDY66P5IvtoVxu
1f5PKinioS7RjgWnuIWyUBmoSG3SpzU1MFnRbo9+pQ1qJw+eNPQtPTj+RyoBwmuAtdUU7i6Be6Oz
UQ/sVoLHBezByYOdTEUOgfocgbNX8v6XJuTXz1Fzrk1AYRvhMdFXmJaS5cvpk3+LW3/8ncy+/j6Q
DAVzDN2I3qp2U5atquBUelKh59HHdHBN/LTxDMB5ISJF5l/fEdfuIdrzr+ZFu2QrIl6T3KFXMceX
qmnmmz1/oLxwE7ft0up+nchVcSiYrgfCaOaTEjnHI8KwQ+9lQGV2pzQpDn94QKDTAWp+UIDEIOaw
cBagHxOS3CR8Nrueo34DLQPcEuoKe13EOO8FdgS3qtXBUB9WqOd84UVGTir+hRcaUg8B2y9dJoTM
nPZW1pTCj9m9GKBQUyQFLMaQO/25t27yWOHCaw40zk2OTh92hLgkFqJcMfBbDhLIgrTTGp35VyO6
vMEGOY9M/8I89FY6Km6izK3s2KJMFpJHA+HrOHtmUoFba28krpN2YKp072LMKK1zVCIHFySfoKDZ
0PmZ8PnL10F7QB3tOqzFkE6I4UF3+jpXROxnKy9SPbqHTgL6W/a1qx1yer69SeHhpnL1FhscBl+N
6ePWnw/0vfsdG+kJ+eEi76OE2GmmufhX1W4GuN1iBtJG2lvY5CIdisjBuYgGU0JKNQnkI90F/Jq6
l/mJYNzAPqKdjqausNPRMEgON0g0ki7NQiDynJjhgZgYmPQtYN1QPKfBl6r+KcZOw7WfkWZJkkKu
WZN9Kw0Txj0Eoe9P3N24MFN3NZkLdzyLVhzn4UbGX5qOCDglVrXm6rCLxkTLnMRs5HAmV93uyBDk
sIs1RT3H7orLCk+IMqtV9KOWP8f6E9IHKGf+lXf09NxcfT8ZHqAYF0l3PyxvGtzDFP4SqrVfJZJU
ECjJ5XczbIG9eSsUuGMx8JE8ZCHJWGsZKx+wAXRZMO7yaV80UfyXQxYQ45hKBKYVq6I/CKN/DTCn
amlsYRFZWNGUGBHOMeEgYkqo1FGWJMEHAn1MjDapYNTXuOknanFL03teouMsUdqdhflfPb/mQ7tW
GhGzqXRX1sH7AlWKB/O36A4MM0NA24E82qyUsuYAUfr0KVi3vG+Ql1+s9kObe7fanNG1tIIQAHyG
rxVrverCpi5IjxY4fFKGDlUm5yVp/O0Nw6Z8sQf7ImrO/BpBjWaYWB/0SEfb0wX2JilFrUHpf/ia
vOPQsHMq/rwHyJDYbnNmmOrUi2s7EE6FZ4gmkfxVunNm8qnKF+OdC+pqKWAACSrtZUVf+YRQj60w
GL/i6Aa1ME2aviVPwDmuDgYoeC73bGbWWmiKB+vh2YPeVuu6yuL6QvQNVMZ933IiVdPL+hnVSNt/
0b5EUyZFxeI+F2X2T5sSRAkLYts2xxpnUG8XZ/vz7edCM8zp8ypXS0+K/y0w8pZgWWSouI+kcf+i
PTpI+lLx97IrLuFprBfYxeyP3gFHxuaG9g8CixwWtldsP0gsUSaZ3MB/llseWVvI+jri9uYTM7Oj
9YAwFwTXpyG5NELIi8VHnsldsccBIWyd4JZslV8f9QpuIihWflYhormBTFofiEl9zmjEHKMq+Xrt
zEYQJGkJc1O6epR+iFTnLqeOSwH5VEev81zaCzFGoTUPotAm2kbAv7ud0fWT5JoRq+WDY9kdl4aF
6eNj5t4x3gmVQ0DO5hwkqe3xQf8i/kvxK4XfcQZUAPhT/pX2rydaURZ+CdtxWf2ubWUPEanhm4Em
S8SudQyLjSnU8gqAB9QbTX6L/fcr1o4BqE4VyGdWGJ8hfat5/T9Suo7ndK19ZL1R8YT4jD0mbJ6A
oyLrS8dXuyYlXE4dZ6IAbcKEIUKXPo88Y6gi+R32aHus6gSG4UMW8aj7rDn5jA3hTcqnvwny+NFo
fHptVAwS8mjm/rnfhrixZbjsVEOYmO0T9fO4HcTBHZqt6nkRvsS0h1jgtGrr6Kfq9GpvAwk1lM+T
xzFC1brN+fTxSVRMXt2nAbUZe/VLfy+x9wVqXqBCMW6LWfiz4MMTosiOSovt+9kqY3q9gjfw95hU
SdxPd77AE+mSnEHHHEjU70g7fUjNC8xK9BAq6LdoDQDSD6F+tVy1OEvZw/vbwrv+Muz57GIqsKZV
A3k1YJDSNfm6s+sQ1PuzomfG1zkPUmXvdNK1+PGSaiXMxzmsjNRnKxEh6ghnoyid/1mcRGlezZs0
2Sw+/MpU+HaaOAdJudG2WHhn+l7Z6+hhBfrLBx4wwNHH5vcwPLVkDW9kN8sN1VF0omaAWvMAJhg9
5v2hNVyGxzSOcvPlWMn+i5TF5E69s7lBfAiKOzPsWFgwV+qeK2ijG9rI6ZMLqHgqhXirVLIYi9uH
dmLxYzH4sZ3LVhxCV+mdvabyMaTnIj8swkIK3L76lUW7w379lSBN1F/f3J8NNM/5U4E+R9y7IZ1A
agceNA3sbXcLJcAXxBp/hcAfMsWgIMx2OZ8PwgdP39p9hn9fOhplFncFIboDHgv0L9Q6wnUg20go
trhoC7HVNxhU6V0QR/Waajl380lcvHlabZJRmge4gTSYOjTWleo35tOo6UG6QEv2q0Is12OYHzaE
kMuGEDz0V2OeQadTEDOQfNVCwflkehRV54Md1fK5ycaRdbaLCidCsYIy1TqJ0StDJG1VjKtWnMjq
IFS7rS5ynIgITJzKWS61nt6Z/Gyrut9zlI2DWagMNpuEcseOW5AByQWYm6l1nt4sjuqWC2LvPUUo
uNxPNquq6NsKNyn/LxoYXW4moCAu2GxSWoAqww8k1qcx6fVoNtEPshemBLx5vGhv9I2YHWXiqSv+
0pqZDH14u+i6kmTFFNH2/wfdgnxvWTlxA9JNsBX93cDN2CPN1gy8wx7dDgrfwTGEsx6UdUQFzLMN
bwMK0zVx+bK4VmpcAED+lgypSLQJmgaYaVmXbUNe4JR1fvmH4+SJx+7+8lfNPiX4neaM99Y8g5s5
oJJkxHw8t2O4aP83UqKZkdU3yCLpQPQv+DWRrTqvc89XDZAjFI38dWMFt06Oaf90cKUvulotnppv
GRq3rFKAcUHKQ2TXzsUdmjqwmxQG+dv7ISlJDwjl3RsN6nCx4E4H5rmfYSaq51vjcDnpZ17PVZgd
E4NXEUlqCtz+1bPNEC/DIuSdCVbALFGggDzO+h5MtmjelYWLAimdB1M//QbtzVY/a6bFdHFQgZFY
PA/gPJUNbY/xiP3TLiRx8EG0saM5go0FAcbFsIHD3XTLpZ+4g444rO7fW8OAJRChuTVAr9EhLstO
YPLMTolc9F0KaqA8PBAAdacyY+cX2tZ9TuxZh0U7ksshDbb47LVFnTP90qpHiYCQqRgYm8FY/pEN
Qv5iiaAvW0JQpxor44PipBhk25XkPiaZid2KitBbP0YwUGy4qEcWJ7QhczzDb4gOmFC7qvjujNJ+
7RenGaRnLdUAvO2aZpVr0SlDs+aQ/UcBFlXAqVrz4XFDHFMheHoMyS5x+xFHbntc8/9HldqYX0kA
u9XUvLW7JY6EeXEAt9lYL336pzISLFN85by64PlVcXLxzA9KXiUI1tIXyt8xyBwdeBi7ZvZp0Abr
U0h2nONuso69iSC35eVRTE8uBjmf55sEDuufGS7xFZ4mJ7VDYINelfsSwWkXRm9LqqECeFZCMk5d
fyPjGSyS3lT8ERnnVPaVshLYxCsly8uqz1morchvbx6J8g6B6PfZ57i4COxs8T3biB/Q6bXK6fyC
4hiMIj7mvj51kDvY38EBDuffs6+hao63eLbKsiA2tJVeO5euoswbcRRENOLVonDViRpyKoUIgILs
7MsZEJS++TvoakrMA8nhwRy80JBPQf0it6ZfmIvcX5Y7AMgWPbdvN8EkzyOx8s0AB7FXq1upn+ix
cnT4YCI5NJUrBb4P0hkpzdRaWj4AjUPrZEQJ6s8jYMcNNHXSnzp6aoDhLdeaaerlLy/CwN+SuWQn
FKv3Fj9OT33Py3xFVg4xczuzJ+b2qIyirkVFxFW3CityL9+iBEIjXv+PP02OGkmlbe4ki9lTPmBL
MXyXkBuaeYrHpPnRNjDuLgtK798fW/BiQFX70ox5qfpVqpZGz23ULnlH7XZ3g4ADVNTtRThHVtIV
lEkp519UF6N37Vvf56wT+Y9JmtvmDEQEza+18kiREB8a4uekvX3ndaM4lV8w9FduF0igQNWATg5y
gvxhkAYi9W/vmRVe25MZQEBC6/cha8QyQcC87qLMechT/kPiM7DXhM9t+s6qlurFeyRFvZrAkZTO
HiPaAGS1zqWFKeyYLDzw5WzsPi6w5UnMxzb6QeksVKKH1Adq3fkbyadHlqI2sb0edf/mNEt5x2ON
8XwoyayWDGyOmuRjQnf30z4yDptclFJQ4CtptM9sCjkq6j0plldt1y3JQq7oObe6ds+d72FPpDGv
ikka18d1TnzvgQ1j828D/qVNd96AV6iTizjebK1P0RDpJzFyZpmPfG607YP0YdWtHO/azi5GUKI+
7v+sYNIXzQkQRFALKKaHmVbBmXTHyfTRKKN2ewdUhuDtiTvr0Gvl8rzfD0y3RIbiPVMGhRn9xvmM
rrAE7FNbkr0AfBFeeXgXS7a1IPZiiKAIH3bWDmJbM59F/66WljF4NOFQ9L0IYzVXrX7Ud3j/CZHQ
ktX7Fu49rITq0H+nEayWAPtG/F8JFuBo1Vm47Q4UMIznDFqBzmFODXkB38DPkpGRjk5kEVSjHX2B
hhxR6MfpzHSfyexZQvXrPHHJa6sGP5hJNgLMBUBxFY7J1XsskvC5q/oKPyl/sbpNBhoWGFFmd7sA
Sv2C6nTM6tZk8Rf7DXqK/MWJmXF5RAODdzWtjCofSDBfi6dm7BRt8+YoO2UfHCZuPwfBaO8YEMKI
ttXbsCjHCmNI2MBHg8OrSWosQIzCg+vz7Bo2jNgjks2Aum4BMX73QoNzPLQgj2H11hhDlrlMl6fD
3SeRjDAiZakgeiK3UgVUI9CkUg3nsS8Ut/rFgho1PPUiBsv6s9JltMavVGtAIQVQm173k7olupwF
YetajCvwNfla0QkxABYEeDTVW8N3UHNlaoET8ghJ3tev7sbfUMtQL7nc91IRJXveeaDeZyhkomPz
0CyhU37UJmePdHY+sBaUQef38gTyc+jrxfT+ioglth7SBWqPri+QhrcLGxQvstaVaZMZg2loSdJy
WX7OZhOkuYJg/cbrs5XSDDMKr+Nl7CjGkOr8aQdCRGCV941Kwmt0yM0o+DaPOlcqC9TKYFH0IMwh
7bQT4YnuV5W6ckzIs+3PMwF7ofxlnPLeIWXFJSKGuxJypyrSiIGYrZw/x+3q81wHiAA5s3cUX7Hv
oQm0RLTdi/xSeZ4GmkJGrdxIwx2imgjE4flouVKUoaUGI1sGdCCx0g99X4y3CPBvvSCylAzn4vQ+
XOyCuxpdXHuIUVIQNPXcGhgtBDcrSx8JAr7onpprLSMg+MdMWoixl8rbP9cX0Hx8fsVpV575us0Q
tM7KNNV/DCcMkPlrc4C2uaubiGepiFEjXUaBUSCOMEEyPfXAUhkfaFbhB+zIDPrAY01lReWe+ItK
6aQpXgc2VZ65Ny1rC8mLhng6BiUSyJ/W1zzRe72rKX0xgf/SxDyhADXJufKeE817UQYh8X3zM93r
bgSpiWfXWuh0Jutq5cdM8b5LTaE/Zqhd00I/pBTCNjTh60Ha+1/Ql63+SfpPHoXm2NtBV1KiWZTE
pjIbPJwl+veVX1HuuNODiobXW0DgIWhsMJi4IpITYzW+UuvVWZTs0nEndv4UXKNG1hRCHMDmhVSq
gLl/bUO+K/3CwD9ZOKCxDLGATcBrjII5RwUpNEpSODZAx7XLSfwsWnGJFjWr6zZrb/iKq4mgHc5+
yUcRAkhVxLtsLMD5fNZGAx+s+FCGd9ctZHvCt97/vTCPtoRIPGyw0cxwexBKmzpH5UO433CwHruM
81riP0Rxzm1s1M8CwxaS+BEVr86Oa+e/hT/Yb9LkMYWr7U5O1stQxPd2foduiG392TVvVmoWU1wB
Cm0pTjwY/hhpgLaoieLYyuQwpM17dw1BRbEuKoeIzVHz/m8ZLqGIGgy+0vKUxJo5O6TgoKAU31hk
6lWoZ0ENOuD5u+J41lDNAEoZc/u3w9MMXRwAWHfOwBeEKDjo2l6vbyNvbJEbAB97RPBjSVUb/NMu
oyoOQC79wOLGAFlZFPprTHxu4zdQ8toggO368qTtfWzUZfqZV8jP5NHUfAEbuMzbpBJ2m6fcoOdm
gwC+stW6Dmq8X/5DL4wKbQktR2iyorfEMid0/wXVZ1iSkQjLed9BvjQg53flhdjQF1priNfX01UU
gwkH0hg//e1AopiWJcRg62NAb4v1lKx/xUw84o/zaUiWM1V24p/wM6dLX5I18+xSfPovuigJkWg9
iynVBwO8gXi9Ul3XOY8a/hgk2pLcwqOQRk75UjWj7np7r7T4GN7echWPkJFWryG6LzXUyvWgeAKl
hDF6sOqgTHVv+iFoG/J7Qd7ClyMr7Ec+zC8u4nTzWBLFjYQDqWirfGuf0QJRGJguZC+4/IUm5hN+
DHnoAZmNaoyOJWHVcBJ5KLQdxhfBv15oUBcSabB+4zFj1SoJTd0fkwW/V5gZCVyKfpvx6PO/Ijip
wUbfzBbkH793LM/3TQMvaRAvwxreUEisY3jdAuDNSF2FcW0af00YVYsw7W46/8nnoyQbYtbrbvoy
tprv59j5JSztPRg3VPvC3n9xn4xsF7v8wo4Oi3Ye9J1dSd06zNctJOSxLJZ+4INKrwL0h0fNVjdv
/xc/BPzjaoVmOvDbsbCxR9XFda8CHorkDrVu2KW8ErcP5cBt3CWVd6a1Mlnbh0oRYvSKEq/k6PRi
qIGllROSP7qypvFowKvXCSW3C1TpJIyRERIBdqk0qrSyCXlFnLoyXtjY4z8OhtWiZ0Jr3IzOjbgt
3qJbGtadJc9HsFj+6v6dJM+WX4DQh9ZwO6OvAUDP2aeOEO34wlDNitDkpo+Sr1J+DRLioWSV7gvd
aCuMqiHrtKWuqCYdf0HLSytzuqYxn6SR628o+o2vLDB6Vs5FiAG5NccmMh1zx9Ss0z/jxGfai0o2
6SpQVkE92HofaN5r1gtz4v42YFYvZDQK9zsyAtsdOKrbuyveix06lkryzmcatnV+9s/JPapzYN01
JRciciCpwfQlbKcj45+iRJKkxYs416HrBoICqx224kM5cvph2etK/DIT+Wwx3E0/vbvXYKmtKZlH
BAHwIFBKOo3/dpChdkAyP2V3Np0XegFCBWu2pvDuys964/+/oj+WDP/gI3NBukKGdAIdSVvyGCTP
8XGFG8fzGsmsd7I5sfWVUSt+bpX4kg0Fu223JHNn0u5Us6kYcrF6gk1xumJKh7QMzZjRYUYuWNc/
NVJJ0mRHbrWcHClA0u7UZH4SON5Osl7H2gJs9vHfnrjnH1ootesb2C9LHOrlyT97KFiDJA7qSrrV
+mRjC/mPOCBCkmo8Ff4NwKYdXDa8J1SKA+E6E+iLPLnaEeNylHWLwLXDV3XwoXs8vRt0D6lu+o1U
ErJfKvkzIPjvJsMmPXYCHV/ggY5uQRgwK8ypEivlV/pFtfz6C+7wfN1M+q15SDiNJygG0dacLcgD
wRKSV2jgg8qmuXhnU+ehbLijLeOD2HZaAc1YvODmhVoImyLnMtltnKo136QZYIajebUOg9PJpcA/
X3k6FrOyNaNuPiLglAYzkST1OBID4RsC2YbUMLPF3oPAIyRiaUAohqImo/FdpGk3Fc3LCb+VHs+O
Ej38ylFILREkHf0wC4kT93JJ+6ZUZrUgVL/WqsikvR9EWlPseUdJYRaMP4dGKX4582CnDhEoOorC
z5Z1KRJf0coyjGUGvv74XlYyckLBZC9DVyXCOLFZ+/Jj+6ii1OQaOsU+HJWHyvzwVOynArZSAcAb
n8OcMWSMptHtrvNw2ayLoiJ/d7SXEnW8OJzl0ntoAL+2h45MV0+A3axvHDZGC+3dIaUb/+LrlZIO
mrTDayN/YTj6x0c8KSG9bcb88JFTVURTKmjrlz7UFD79eLH50gilGhYWOcHUo2b0yGIiC3dD44oM
527OPyvQLIE4HjjgtrdYB8EpYO8OBJ1Y6pWT6Izbg3J6iMhHIp7kNCdv7DyjYcJ9PsGup4QdT+3u
eVkNYGs38Vukxkc51y7iF8CPUugm3+1EDNdvFpcIgqZP8H32fPTp8tT92mdvd4KVkXtoxXy71bc=
`pragma protect end_protected
